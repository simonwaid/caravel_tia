magic
tech sky130A
magscale 1 2
timestamp 1646925174
<< metal1 >>
rect -7840 11160 -7830 11400
rect -7550 11160 -7140 11400
<< via1 >>
rect -7830 11160 -7550 11400
<< metal2 >>
rect -3800 13260 -3650 13270
rect -3800 13080 -3650 13090
rect 6220 12150 15900 12160
rect 6220 11980 6230 12150
rect 6380 12130 15900 12150
rect 6380 12000 16070 12130
rect 6380 11980 15900 12000
rect 6220 11970 15900 11980
rect -7830 11400 -7550 11410
rect -7830 11150 -7550 11160
rect 16000 10970 16060 11040
rect 15350 10960 16210 10970
rect 15350 10750 15360 10960
rect 15610 10750 16210 10960
rect 15350 10740 16210 10750
rect 16500 8630 16640 8640
rect 16640 8470 17200 8630
rect 16500 8460 16640 8470
rect 11920 -4010 13810 -3990
rect 11920 -4330 13480 -4010
rect 13790 -4330 13810 -4010
rect 11920 -4350 13810 -4330
rect -6740 -4500 -6160 -4490
rect -6740 -4600 -6730 -4500
rect -6610 -4600 -6160 -4500
rect -6740 -4610 -6160 -4600
rect -22080 -7390 -20410 -7380
rect -21850 -7650 -20640 -7390
rect -22080 -7660 -20410 -7650
rect 9690 -7620 10490 -7550
rect 9690 -7910 10240 -7620
rect 10470 -7910 10490 -7620
rect 9690 -7950 10490 -7910
rect -21500 -13730 -21360 -12950
rect -20150 -13730 -20010 -12930
rect -18800 -13730 -18660 -12950
rect -17450 -13730 -17310 -12930
rect -16100 -13730 -15960 -12990
rect -14750 -13730 -14610 -12990
rect -13400 -13380 -13260 -13010
rect -13400 -13510 -13390 -13380
rect -13270 -13510 -13260 -13380
rect -13400 -13520 -13260 -13510
rect -12050 -13400 -11910 -13010
rect -10700 -13060 -10560 -12850
rect -11210 -13070 -10560 -13060
rect -10960 -13210 -10560 -13070
rect -11210 -13220 -10560 -13210
rect -12050 -13520 -11910 -13510
<< via2 >>
rect -3800 13090 -3650 13260
rect 6230 11980 6380 12150
rect -7830 11160 -7550 11400
rect 15360 10750 15610 10960
rect 16500 8470 16640 8630
rect 13480 -4330 13790 -4010
rect -6730 -4600 -6610 -4500
rect -22080 -7650 -21850 -7390
rect -20640 -7650 -20410 -7390
rect 10240 -7910 10470 -7620
rect -13390 -13510 -13270 -13380
rect -11210 -13210 -10960 -13070
rect -12050 -13510 -11910 -13400
<< metal3 >>
rect -3810 13260 -3640 13265
rect -3810 13090 -3800 13260
rect -3650 13090 -3640 13260
rect -3810 13085 -3640 13090
rect -3800 11920 -3650 13085
rect -270 12160 -30 12170
rect -270 12150 6390 12160
rect -270 11980 6230 12150
rect 6380 11980 6390 12150
rect -270 11970 6390 11980
rect -270 11920 -30 11970
rect -3800 11710 -30 11920
rect -3800 11700 -230 11710
rect -7840 11400 -7540 11405
rect -7840 11160 -7830 11400
rect -7550 11160 -7540 11400
rect -7840 11155 -7540 11160
rect -120 10960 15620 10970
rect -120 10750 15360 10960
rect 15610 10750 15620 10960
rect -120 10740 15620 10750
rect -120 7670 310 10740
rect -4200 7530 310 7670
rect 13470 8630 16820 8660
rect 13470 8470 16500 8630
rect 16640 8470 16820 8630
rect 13470 8390 16820 8470
rect 1770 4330 2020 4340
rect -310 4170 2020 4330
rect 1000 2580 1620 2660
rect -12120 530 -6490 540
rect 1520 530 1620 2580
rect -12120 330 1620 530
rect 1770 720 2020 4170
rect 1770 520 12780 720
rect -12120 320 -6490 330
rect -22090 -7390 -21840 -7385
rect -36360 -7650 -22080 -7390
rect -21850 -7650 -21840 -7390
rect -22090 -7655 -21840 -7650
rect -21620 -8530 -20990 -6340
rect -12120 -7380 -11840 320
rect -9410 -4500 -6600 -4490
rect -9410 -4600 -6730 -4500
rect -6610 -4600 -6600 -4500
rect -9410 -4610 -6600 -4600
rect -20640 -7385 -11830 -7380
rect -20650 -7390 -11830 -7385
rect -20650 -7650 -20640 -7390
rect -20410 -7650 -11830 -7390
rect -20650 -7655 -20400 -7650
rect -21620 -8790 -10960 -8530
rect -18620 -9560 -18610 -9140
rect -17930 -9560 -17920 -9140
rect -11210 -13065 -10960 -8790
rect -11220 -13070 -10950 -13065
rect -11220 -13210 -11210 -13070
rect -10960 -13210 -10950 -13070
rect -11220 -13215 -10950 -13210
rect -36660 -13370 -20670 -13350
rect -36660 -13380 -13260 -13370
rect -36660 -13510 -13390 -13380
rect -13270 -13510 -13260 -13380
rect -36660 -13520 -13260 -13510
rect -12060 -13400 -11900 -13395
rect -9410 -13400 -9080 -4610
rect 12520 -7610 12780 520
rect 13470 -4010 13810 8390
rect 13470 -4330 13480 -4010
rect 13790 -4330 13810 -4010
rect 13470 -4335 13800 -4330
rect 10230 -7620 12780 -7610
rect 10230 -7910 10240 -7620
rect 10470 -7910 12780 -7620
rect 10230 -7920 12780 -7910
rect -12060 -13510 -12050 -13400
rect -11910 -13510 -9080 -13400
rect -12060 -13515 -11900 -13510
rect -36660 -13530 -20670 -13520
rect -36660 -13540 -25550 -13530
<< via3 >>
rect -7830 11160 -7550 11400
rect -18610 -9560 -17930 -9140
<< metal4 >>
rect -10180 16050 -9260 16070
rect -36230 15010 -9260 16050
rect -10180 11940 -9260 15010
rect -10180 11400 -7540 11940
rect -10180 11160 -7830 11400
rect -7550 11160 -7540 11400
rect -10180 11150 -7540 11160
rect 5830 2800 8110 2840
rect 5830 2110 7210 2800
rect 8070 2110 8110 2800
rect 5830 2070 8110 2110
rect -12110 -1770 -6080 -1750
rect -11810 -2780 -6080 -1770
rect -12110 -2790 -6080 -2780
rect -18611 -9140 -17929 -9139
rect -18611 -9560 -18610 -9140
rect -17930 -9560 -17929 -9140
rect -18611 -9561 -17929 -9560
<< via4 >>
rect 7210 2110 8070 2800
rect -12610 -2780 -11810 -1770
rect -18610 -9560 -17930 -9140
<< metal5 >>
rect -36460 16840 93590 19280
rect -12640 -1770 -11780 16840
rect 3720 13820 4440 16840
rect 6990 15680 8180 16840
rect 35360 15160 36180 16840
rect 49920 15080 50740 16840
rect 64330 15240 65150 16840
rect 78370 15180 79190 16840
rect 92550 15360 93370 16840
rect 7186 2800 8094 2824
rect 7186 2110 7210 2800
rect 8070 2110 8094 2800
rect 7186 2086 8094 2110
rect -12640 -2780 -12610 -1770
rect -11810 -2780 -11780 -1770
rect -20580 -13776 -19740 -6270
rect -19370 -6890 -18570 -6390
rect -12640 -6890 -11780 -2780
rect -19370 -7700 -11780 -6890
rect -18610 -9116 -17930 -7700
rect -18634 -9140 -17906 -9116
rect -18634 -9560 -18610 -9140
rect -17930 -9560 -17906 -9140
rect -18634 -9584 -17906 -9560
rect -8800 -12450 -6100 -12020
rect -20580 -14374 -19376 -13776
rect -20580 -16740 -19740 -14374
rect -8800 -16740 -7620 -12450
rect 14490 -16740 15950 1420
rect 86310 -16740 88850 1170
rect -36770 -19180 93280 -16740
use cmirror_channel  cmirror_channel_0 ~/code/caravel_tia/mag/currm
timestamp 1646921651
transform 1 0 -7150 0 1 -4140
box -60 -11100 19842 4124
use eigth_mirror  eigth_mirror_0 ~/code/caravel_tia/mag/currm
timestamp 1646921651
transform -1 0 -10420 0 -1 -9430
box 10 0 12180 3580
use isource  isource_0 ~/code/caravel_tia/mag/isource
timestamp 1646921651
transform 1 0 -36170 0 1 -1620
box -280 -4830 23120 15920
use outd  outd_0 ~/code/caravel_tia/mag/outd
timestamp 1646921651
transform 1 0 37150 0 1 700
box -30220 -60 57040 15224
use tia_core  tia_core_0 ~/code/caravel_tia/mag/tia
timestamp 1646921651
transform 1 0 -5400 0 1 12420
box -1860 -11680 11730 2790
<< labels >>
rlabel metal3 -36650 -13530 -36380 -13360 1 I_ref_out
rlabel metal5 -36510 -18610 -35610 -17020 1 VN
rlabel metal5 -36200 17300 -35300 18890 1 VP
rlabel metal3 -36350 -7640 -35860 -7410 1 Dis_TIA
rlabel metal4 -36170 15070 -35340 15970 1 TIA_in
<< end >>
