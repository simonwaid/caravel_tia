magic
tech sky130A
magscale 1 2
timestamp 1645630008
<< nwell >>
rect -812 -1137 812 1137
<< pmos >>
rect -616 118 -416 918
rect -358 118 -158 918
rect -100 118 100 918
rect 158 118 358 918
rect 416 118 616 918
rect -616 -918 -416 -118
rect -358 -918 -158 -118
rect -100 -918 100 -118
rect 158 -918 358 -118
rect 416 -918 616 -118
<< pdiff >>
rect -674 906 -616 918
rect -674 130 -662 906
rect -628 130 -616 906
rect -674 118 -616 130
rect -416 906 -358 918
rect -416 130 -404 906
rect -370 130 -358 906
rect -416 118 -358 130
rect -158 906 -100 918
rect -158 130 -146 906
rect -112 130 -100 906
rect -158 118 -100 130
rect 100 906 158 918
rect 100 130 112 906
rect 146 130 158 906
rect 100 118 158 130
rect 358 906 416 918
rect 358 130 370 906
rect 404 130 416 906
rect 358 118 416 130
rect 616 906 674 918
rect 616 130 628 906
rect 662 130 674 906
rect 616 118 674 130
rect -674 -130 -616 -118
rect -674 -906 -662 -130
rect -628 -906 -616 -130
rect -674 -918 -616 -906
rect -416 -130 -358 -118
rect -416 -906 -404 -130
rect -370 -906 -358 -130
rect -416 -918 -358 -906
rect -158 -130 -100 -118
rect -158 -906 -146 -130
rect -112 -906 -100 -130
rect -158 -918 -100 -906
rect 100 -130 158 -118
rect 100 -906 112 -130
rect 146 -906 158 -130
rect 100 -918 158 -906
rect 358 -130 416 -118
rect 358 -906 370 -130
rect 404 -906 416 -130
rect 358 -918 416 -906
rect 616 -130 674 -118
rect 616 -906 628 -130
rect 662 -906 674 -130
rect 616 -918 674 -906
<< pdiffc >>
rect -662 130 -628 906
rect -404 130 -370 906
rect -146 130 -112 906
rect 112 130 146 906
rect 370 130 404 906
rect 628 130 662 906
rect -662 -906 -628 -130
rect -404 -906 -370 -130
rect -146 -906 -112 -130
rect 112 -906 146 -130
rect 370 -906 404 -130
rect 628 -906 662 -130
<< nsubdiff >>
rect -776 1067 -680 1101
rect 680 1067 776 1101
rect -776 1005 -742 1067
rect 742 1005 776 1067
rect -776 -1067 -742 -1005
rect 742 -1067 776 -1005
rect -776 -1101 -680 -1067
rect 680 -1101 776 -1067
<< nsubdiffcont >>
rect -680 1067 680 1101
rect -776 -1005 -742 1005
rect 742 -1005 776 1005
rect -680 -1101 680 -1067
<< poly >>
rect -616 999 -416 1015
rect -616 965 -600 999
rect -432 965 -416 999
rect -616 918 -416 965
rect -358 999 -158 1015
rect -358 965 -342 999
rect -174 965 -158 999
rect -358 918 -158 965
rect -100 999 100 1015
rect -100 965 -84 999
rect 84 965 100 999
rect -100 918 100 965
rect 158 999 358 1015
rect 158 965 174 999
rect 342 965 358 999
rect 158 918 358 965
rect 416 999 616 1015
rect 416 965 432 999
rect 600 965 616 999
rect 416 918 616 965
rect -616 71 -416 118
rect -616 37 -600 71
rect -432 37 -416 71
rect -616 21 -416 37
rect -358 71 -158 118
rect -358 37 -342 71
rect -174 37 -158 71
rect -358 21 -158 37
rect -100 71 100 118
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect 158 71 358 118
rect 158 37 174 71
rect 342 37 358 71
rect 158 21 358 37
rect 416 71 616 118
rect 416 37 432 71
rect 600 37 616 71
rect 416 21 616 37
rect -616 -37 -416 -21
rect -616 -71 -600 -37
rect -432 -71 -416 -37
rect -616 -118 -416 -71
rect -358 -37 -158 -21
rect -358 -71 -342 -37
rect -174 -71 -158 -37
rect -358 -118 -158 -71
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -118 100 -71
rect 158 -37 358 -21
rect 158 -71 174 -37
rect 342 -71 358 -37
rect 158 -118 358 -71
rect 416 -37 616 -21
rect 416 -71 432 -37
rect 600 -71 616 -37
rect 416 -118 616 -71
rect -616 -965 -416 -918
rect -616 -999 -600 -965
rect -432 -999 -416 -965
rect -616 -1015 -416 -999
rect -358 -965 -158 -918
rect -358 -999 -342 -965
rect -174 -999 -158 -965
rect -358 -1015 -158 -999
rect -100 -965 100 -918
rect -100 -999 -84 -965
rect 84 -999 100 -965
rect -100 -1015 100 -999
rect 158 -965 358 -918
rect 158 -999 174 -965
rect 342 -999 358 -965
rect 158 -1015 358 -999
rect 416 -965 616 -918
rect 416 -999 432 -965
rect 600 -999 616 -965
rect 416 -1015 616 -999
<< polycont >>
rect -600 965 -432 999
rect -342 965 -174 999
rect -84 965 84 999
rect 174 965 342 999
rect 432 965 600 999
rect -600 37 -432 71
rect -342 37 -174 71
rect -84 37 84 71
rect 174 37 342 71
rect 432 37 600 71
rect -600 -71 -432 -37
rect -342 -71 -174 -37
rect -84 -71 84 -37
rect 174 -71 342 -37
rect 432 -71 600 -37
rect -600 -999 -432 -965
rect -342 -999 -174 -965
rect -84 -999 84 -965
rect 174 -999 342 -965
rect 432 -999 600 -965
<< locali >>
rect -776 1067 -680 1101
rect 680 1067 776 1101
rect -776 1005 -742 1067
rect 742 1005 776 1067
rect -616 965 -600 999
rect -432 965 -416 999
rect -358 965 -342 999
rect -174 965 -158 999
rect -100 965 -84 999
rect 84 965 100 999
rect 158 965 174 999
rect 342 965 358 999
rect 416 965 432 999
rect 600 965 616 999
rect -662 906 -628 922
rect -662 114 -628 130
rect -404 906 -370 922
rect -404 114 -370 130
rect -146 906 -112 922
rect -146 114 -112 130
rect 112 906 146 922
rect 112 114 146 130
rect 370 906 404 922
rect 370 114 404 130
rect 628 906 662 922
rect 628 114 662 130
rect -616 37 -600 71
rect -432 37 -416 71
rect -358 37 -342 71
rect -174 37 -158 71
rect -100 37 -84 71
rect 84 37 100 71
rect 158 37 174 71
rect 342 37 358 71
rect 416 37 432 71
rect 600 37 616 71
rect -616 -71 -600 -37
rect -432 -71 -416 -37
rect -358 -71 -342 -37
rect -174 -71 -158 -37
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect 158 -71 174 -37
rect 342 -71 358 -37
rect 416 -71 432 -37
rect 600 -71 616 -37
rect -662 -130 -628 -114
rect -662 -922 -628 -906
rect -404 -130 -370 -114
rect -404 -922 -370 -906
rect -146 -130 -112 -114
rect -146 -922 -112 -906
rect 112 -130 146 -114
rect 112 -922 146 -906
rect 370 -130 404 -114
rect 370 -922 404 -906
rect 628 -130 662 -114
rect 628 -922 662 -906
rect -616 -999 -600 -965
rect -432 -999 -416 -965
rect -358 -999 -342 -965
rect -174 -999 -158 -965
rect -100 -999 -84 -965
rect 84 -999 100 -965
rect 158 -999 174 -965
rect 342 -999 358 -965
rect 416 -999 432 -965
rect 600 -999 616 -965
rect -776 -1067 -742 -1005
rect 742 -1067 776 -1005
rect -776 -1101 -680 -1067
rect 680 -1101 776 -1067
<< viali >>
rect -600 965 -432 999
rect -342 965 -174 999
rect -84 965 84 999
rect 174 965 342 999
rect 432 965 600 999
rect -662 130 -628 906
rect -404 130 -370 906
rect -146 130 -112 906
rect 112 130 146 906
rect 370 130 404 906
rect 628 130 662 906
rect -600 37 -432 71
rect -342 37 -174 71
rect -84 37 84 71
rect 174 37 342 71
rect 432 37 600 71
rect -600 -71 -432 -37
rect -342 -71 -174 -37
rect -84 -71 84 -37
rect 174 -71 342 -37
rect 432 -71 600 -37
rect -662 -906 -628 -130
rect -404 -906 -370 -130
rect -146 -906 -112 -130
rect 112 -906 146 -130
rect 370 -906 404 -130
rect 628 -906 662 -130
rect -600 -999 -432 -965
rect -342 -999 -174 -965
rect -84 -999 84 -965
rect 174 -999 342 -965
rect 432 -999 600 -965
<< metal1 >>
rect -612 999 -420 1005
rect -612 965 -600 999
rect -432 965 -420 999
rect -612 959 -420 965
rect -354 999 -162 1005
rect -354 965 -342 999
rect -174 965 -162 999
rect -354 959 -162 965
rect -96 999 96 1005
rect -96 965 -84 999
rect 84 965 96 999
rect -96 959 96 965
rect 162 999 354 1005
rect 162 965 174 999
rect 342 965 354 999
rect 162 959 354 965
rect 420 999 612 1005
rect 420 965 432 999
rect 600 965 612 999
rect 420 959 612 965
rect -668 906 -622 918
rect -668 130 -662 906
rect -628 130 -622 906
rect -668 118 -622 130
rect -410 906 -364 918
rect -410 130 -404 906
rect -370 130 -364 906
rect -410 118 -364 130
rect -152 906 -106 918
rect -152 130 -146 906
rect -112 130 -106 906
rect -152 118 -106 130
rect 106 906 152 918
rect 106 130 112 906
rect 146 130 152 906
rect 106 118 152 130
rect 364 906 410 918
rect 364 130 370 906
rect 404 130 410 906
rect 364 118 410 130
rect 622 906 668 918
rect 622 130 628 906
rect 662 130 668 906
rect 622 118 668 130
rect -612 71 -420 77
rect -612 37 -600 71
rect -432 37 -420 71
rect -612 31 -420 37
rect -354 71 -162 77
rect -354 37 -342 71
rect -174 37 -162 71
rect -354 31 -162 37
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect 162 71 354 77
rect 162 37 174 71
rect 342 37 354 71
rect 162 31 354 37
rect 420 71 612 77
rect 420 37 432 71
rect 600 37 612 71
rect 420 31 612 37
rect -612 -37 -420 -31
rect -612 -71 -600 -37
rect -432 -71 -420 -37
rect -612 -77 -420 -71
rect -354 -37 -162 -31
rect -354 -71 -342 -37
rect -174 -71 -162 -37
rect -354 -77 -162 -71
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect 162 -37 354 -31
rect 162 -71 174 -37
rect 342 -71 354 -37
rect 162 -77 354 -71
rect 420 -37 612 -31
rect 420 -71 432 -37
rect 600 -71 612 -37
rect 420 -77 612 -71
rect -668 -130 -622 -118
rect -668 -906 -662 -130
rect -628 -906 -622 -130
rect -668 -918 -622 -906
rect -410 -130 -364 -118
rect -410 -906 -404 -130
rect -370 -906 -364 -130
rect -410 -918 -364 -906
rect -152 -130 -106 -118
rect -152 -906 -146 -130
rect -112 -906 -106 -130
rect -152 -918 -106 -906
rect 106 -130 152 -118
rect 106 -906 112 -130
rect 146 -906 152 -130
rect 106 -918 152 -906
rect 364 -130 410 -118
rect 364 -906 370 -130
rect 404 -906 410 -130
rect 364 -918 410 -906
rect 622 -130 668 -118
rect 622 -906 628 -130
rect 662 -906 668 -130
rect 622 -918 668 -906
rect -612 -965 -420 -959
rect -612 -999 -600 -965
rect -432 -999 -420 -965
rect -612 -1005 -420 -999
rect -354 -965 -162 -959
rect -354 -999 -342 -965
rect -174 -999 -162 -965
rect -354 -1005 -162 -999
rect -96 -965 96 -959
rect -96 -999 -84 -965
rect 84 -999 96 -965
rect -96 -1005 96 -999
rect 162 -965 354 -959
rect 162 -999 174 -965
rect 342 -999 354 -965
rect 162 -1005 354 -999
rect 420 -965 612 -959
rect 420 -999 432 -965
rect 600 -999 612 -965
rect 420 -1005 612 -999
<< properties >>
string FIXED_BBOX -759 -1084 759 1084
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4 l 1 m 2 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
