* SPICE3 file created from user_analog_project_wrapper_flat.ext - technology: sky130A

X0 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.47712e+15p ps=1.9251e+10u w=2e+06u l=500000u
X1 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7 mpw5_submission_0/tia_core_0/VM5D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 io_analog[3] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.324e+13p ps=1.0124e+08u w=2e+06u l=150000u
X8 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.2544e+14p ps=8.9344e+08u w=2e+06u l=150000u
X13 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X16 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X17 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=1.2544e+14p pd=8.9344e+08u as=0p ps=0u w=2e+06u l=150000u
X18 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X19 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X20 mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X21 mpw5_submission_1/eigth_mirror_0/I_out_1 mpw5_submission_1/eigth_mirror_0/I_In a_192870_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X22 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X23 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X24 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X25 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X26 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=1.2544e+14p pd=8.9344e+08u as=0p ps=0u w=2e+06u l=150000u
X27 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X28 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X29 a_203650_645683# a_201520_649146# mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X30 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X31 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X32 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X33 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X34 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=6.5714e+14p pd=5.12824e+09u as=0p ps=0u w=2e+06u l=1e+06u
X35 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X36 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X37 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X38 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X39 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X40 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X41 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X42 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X43 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/InputRef mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X44 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D0 vssd1 io_analog[7] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X45 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X46 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X47 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X48 io_analog[3] mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/tia_core_0/Out_2 io_analog[3] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X49 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X50 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X51 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X52 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X53 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X54 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X55 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X56 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X57 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X58 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X59 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X60 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X61 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X62 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X63 mpw5_submission_0/tia_core_0/Out_2 mpw5_submission_0/outd_0/InputSignal io_analog[3] io_analog[3] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X64 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D1 io_analog[7] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X65 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X66 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X67 vssd1 mpw5_submission_0/cmirror_channel_0/I_in_channel sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X68 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X69 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X70 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X71 mpw5_submission_1/tia_core_0/VM31D mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X72 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X73 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X74 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X75 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X76 mpw5_submission_1/isource_0/VM12G mpw5_submission_1/isource_0/VM14D vccd1 mpw5_submission_1/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.60134e+15p ps=1.3951e+10u w=4e+06u l=150000u
X77 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X78 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X79 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X80 a_203650_645683# a_201520_649146# mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X81 io_analog[5] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X82 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X83 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X84 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X85 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X86 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X87 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X88 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X89 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X90 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X91 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X92 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X93 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM31D mpw5_submission_1/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X94 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X95 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X96 a_194220_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X97 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X98 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X99 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X100 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X101 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X102 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X103 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X104 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X105 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X106 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D2 vssd1 io_analog[1] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X107 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X108 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X109 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X110 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X111 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X112 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X113 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X114 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X115 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X116 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X117 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X118 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X119 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X120 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X121 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X122 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X123 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X124 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X125 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X126 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D3 io_analog[2] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X127 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X128 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X129 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X130 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X131 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X132 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X133 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X134 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X135 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X136 mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X137 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X138 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X139 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X140 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X141 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X142 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X143 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X144 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=1.2544e+14p pd=8.9344e+08u as=0p ps=0u w=2e+06u l=150000u
X145 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X146 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X147 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X148 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X149 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X150 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X151 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X152 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X153 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X154 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X155 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X156 vccd1 io_analog[0] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X157 a_192870_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X158 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X159 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X160 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X161 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X162 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X163 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X164 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X165 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X166 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X167 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X168 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X169 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X170 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X171 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X172 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X173 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X174 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X175 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X176 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X177 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X178 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X179 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X180 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X181 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X182 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X183 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X184 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X185 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X186 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X187 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X188 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X189 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X190 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X191 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X192 io_analog[6] mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM5D vssd1 sky130_fd_pr__nfet_01v8 ad=1.324e+13p pd=1.0124e+08u as=0p ps=0u w=2e+06u l=150000u
X193 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X194 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X195 a_191520_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X196 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X197 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X198 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X199 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X200 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X201 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X202 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_657119# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X203 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X204 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X205 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X206 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X207 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X208 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X209 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X210 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X211 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X212 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X213 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X214 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X215 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X216 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X217 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/Disable_TIA vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X218 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X219 a_430136_657119# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X220 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X221 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X222 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X223 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X224 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X225 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X226 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X227 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X228 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X229 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X230 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X231 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X232 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X233 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X234 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X235 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X236 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_427670_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X237 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X238 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X239 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X240 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X241 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X242 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X243 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X244 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X245 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X246 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X247 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X248 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X249 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X250 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_192870_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X251 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X252 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X253 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X254 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X255 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X256 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X257 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X258 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X259 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X260 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X261 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X262 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X263 a_189936_651879# mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM14D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X264 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X265 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X266 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X267 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X268 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X269 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X270 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X271 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X272 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X273 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X274 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X275 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X276 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X277 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X278 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X279 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X280 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X281 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X282 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X283 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X284 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X285 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X286 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X287 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X288 a_430136_657119# mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM9D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X289 a_430136_648079# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X290 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D4 io_analog[8] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X291 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X292 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X293 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_429020_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X294 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X295 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X296 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_426320_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X297 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X298 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM31D mpw5_submission_1/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X299 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X300 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X301 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X302 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X303 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X304 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X305 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X306 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_429020_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X307 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X308 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X309 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X310 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X311 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X312 vccd1 mpw5_submission_1/isource_0/VM14D mpw5_submission_1/isource_0/VM12G mpw5_submission_1/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X313 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X314 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X315 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X316 vssd1 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X317 mpw5_submission_1/tia_core_0/VM31D mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X318 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X319 vssd1 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X320 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X321 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X322 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X323 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X324 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X325 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X326 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X327 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X328 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X329 mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/InputRef mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X330 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X331 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X332 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X333 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X334 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X335 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X336 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X337 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X338 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X339 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X340 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X341 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X342 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X343 vssd1 mpw5_submission_0/cmirror_channel_0/I_in_channel sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X344 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X345 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X346 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X347 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X348 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X349 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X350 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X351 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X352 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X353 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X354 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X355 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X356 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X357 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X358 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X359 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X360 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X361 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D5 io_analog[1] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X362 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X363 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X364 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X365 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X366 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X367 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X368 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
D6 io_analog[3] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X369 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X370 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X371 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X372 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X373 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X374 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X375 a_189936_651879# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X376 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X377 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X378 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X379 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X380 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X381 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM31D mpw5_submission_1/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X382 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X383 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X384 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X385 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X386 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X387 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X388 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X389 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X390 a_195570_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X391 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X392 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X393 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X394 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X395 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X396 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X397 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X398 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X399 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X400 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X401 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X402 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X403 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X404 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X405 mpw5_submission_0/tia_core_0/VM31D mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X406 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X407 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X408 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X409 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X410 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X411 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X412 a_430136_648079# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X413 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X414 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X415 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X416 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X417 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X418 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X419 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X420 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X421 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X422 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X423 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X424 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X425 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X426 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X427 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X428 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X429 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X430 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X431 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X432 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X433 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X434 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X435 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X436 a_194220_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X437 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X438 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X439 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X440 io_analog[5] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X441 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X442 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X443 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X444 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X445 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X446 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X447 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X448 mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/InputRef mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D7 vssd1 io_analog[2] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X449 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X450 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X451 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X452 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X453 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X454 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
D8 vssd1 io_analog[3] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X455 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X456 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X457 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X458 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X459 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X460 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X461 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X462 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X463 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X464 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X465 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X466 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X467 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X468 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X469 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X470 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X471 mpw5_submission_0/isource_0/VM22D a_411216_644902# mpw5_submission_0/isource_0/VM3D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X472 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X473 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X474 a_430136_648079# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X475 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X476 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X477 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X478 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X479 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X480 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X481 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X482 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X483 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X484 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X485 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X486 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X487 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X488 mpw5_submission_0/tia_core_0/VM31D mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X489 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X490 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X491 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X492 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X493 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X494 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X495 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X496 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X497 a_190170_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X498 a_188820_640623# mpw5_submission_1/eigth_mirror_0/I_In mpw5_submission_1/eigth_mirror_0/I_out_4 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X499 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X500 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X501 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X502 a_427116_648806# a_426586_651238# vssd1 sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X503 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X504 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X505 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X506 a_429020_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X507 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X508 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X509 a_443570_645443# a_441720_645346# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X510 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X511 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X512 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X513 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X514 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X515 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_187470_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X516 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X517 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X518 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X519 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X520 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X521 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X522 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X523 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X524 vccd1 vssd1 mpw5_submission_0/tia_core_0/Out_2 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X525 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X526 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X527 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X528 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X529 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X530 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X531 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X532 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X533 a_430136_648079# mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM14D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X534 vssd1 mpw5_submission_0/cmirror_channel_0/I_in_channel a_440818_643680# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X535 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X536 a_411216_644902# mpw5_submission_0/isource_0/VM22D mpw5_submission_0/eigth_mirror_0/I_In vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X537 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X538 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X539 io_analog[4] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X540 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X541 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X542 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X543 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X544 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X545 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X546 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X547 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X548 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X549 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X550 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X551 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X552 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X553 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X554 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X555 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X556 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X557 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X558 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X559 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X560 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X561 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_186120_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X562 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X563 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X564 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X565 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X566 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X567 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X568 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X569 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X570 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X571 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X572 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X573 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X574 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X575 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X576 mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X577 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X578 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X579 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X580 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X581 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X582 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X583 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X584 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X585 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_660919# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X586 a_442498_643680# mpw5_submission_0/cmirror_channel_0/I_in_channel vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X587 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X588 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X589 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X590 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X591 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_431720_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X592 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X593 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X594 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X595 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X596 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X597 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X598 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X599 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X600 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X601 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X602 a_201520_649146# a_201520_649146# a_201720_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X603 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X604 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X605 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_184770_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X606 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X607 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X608 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X609 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X610 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X611 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X612 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X613 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X614 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X615 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X616 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X617 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X618 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X619 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X620 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X621 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X622 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X623 vccd1 vssd1 mpw5_submission_0/tia_core_0/VM31D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X624 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X625 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X626 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X627 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X628 a_435770_636823# mpw5_submission_0/eigth_mirror_0/I_In mpw5_submission_0/eigth_mirror_0/I_In vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X629 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X630 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X631 vccd1 vssd1 mpw5_submission_1/tia_core_0/VM31D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X632 a_171016_648702# mpw5_submission_1/isource_0/VM22D mpw5_submission_1/eigth_mirror_0/I_In vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X633 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X634 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X635 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X636 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X637 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X638 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X639 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X640 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X641 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X642 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X643 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X644 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X645 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X646 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X647 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X648 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X649 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X650 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X651 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X652 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X653 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X654 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X655 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X656 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X657 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X658 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X659 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X660 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X661 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_186120_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X662 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X663 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X664 a_443850_641883# a_441720_645346# mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X665 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X666 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X667 io_analog[6] mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/tia_core_0/Out_2 io_analog[6] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X668 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X669 mpw5_submission_0/isource_0/VM3D a_411216_644902# mpw5_submission_0/isource_0/VM22D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X670 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X671 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X672 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X673 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X674 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X675 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X676 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X677 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X678 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_424970_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X679 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X680 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X681 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X682 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X683 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X684 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X685 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X686 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X687 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X688 a_189936_649609# mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM22D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X689 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X690 vccd1 io_analog[5] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X691 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X692 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X693 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X694 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X695 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X696 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X697 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X698 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X699 a_189936_651879# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X700 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X701 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X702 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X703 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X704 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X705 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X706 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X707 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X708 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X709 a_181958_664870# mpw5_submission_1/isource_0/VM11D vssd1 vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X710 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X711 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM31D mpw5_submission_0/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X712 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X713 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X714 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X715 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X716 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X717 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X718 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X719 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X720 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X721 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X722 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X723 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X724 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X725 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X726 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X727 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X728 a_187470_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X729 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X730 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X731 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X732 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X733 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X734 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X735 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X736 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X737 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X738 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X739 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X740 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X741 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X742 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X743 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X744 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X745 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X746 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X747 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X748 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X749 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X750 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X751 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X752 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X753 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X754 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X755 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X756 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X757 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X758 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X759 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X760 a_441920_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X761 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X762 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X763 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X764 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X765 a_203370_649243# a_201520_649146# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X766 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X767 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X768 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X769 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X770 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X771 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X772 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X773 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X774 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X775 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X776 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X777 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X778 vssd1 mpw5_submission_0/cmirror_channel_0/I_in_channel a_441658_643680# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X779 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X780 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X781 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X782 mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/InputRef mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X783 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X784 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X785 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X786 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X787 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X788 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X789 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X790 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X791 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X792 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_645809# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X793 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X794 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X795 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X796 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X797 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X798 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X799 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X800 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X801 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X802 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X803 a_430136_645809# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X804 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X805 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X806 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X807 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X808 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X809 mpw5_submission_0/tia_core_0/Out_2 mpw5_submission_0/outd_0/InputSignal io_analog[3] io_analog[3] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X810 a_435770_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X811 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X812 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X813 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X814 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X815 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X816 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X817 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X818 a_430136_648079# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X819 a_188820_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X820 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X821 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X822 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X823 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X824 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X825 a_200618_647480# mpw5_submission_1/cmirror_channel_0/I_in_channel mpw5_submission_1/cmirror_channel_0/I_in_channel vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
D9 vssd1 io_analog[8] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X826 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X827 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X828 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X829 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X830 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X831 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X832 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X833 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X834 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X835 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X836 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X837 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X838 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X839 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X840 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X841 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X842 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X843 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X844 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X845 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X846 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X847 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X848 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X849 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X850 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X851 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X852 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X853 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X854 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X855 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X856 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X857 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X858 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X859 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D10 vssd1 io_analog[3] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X860 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X861 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X862 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X863 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X864 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X865 vccd1 a_201520_649146# a_201720_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X866 a_434420_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X867 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X868 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D11 io_analog[1] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X869 vccd1 io_analog[4] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X870 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X871 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X872 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X873 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X874 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X875 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X876 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X877 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X878 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X879 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X880 a_430136_645809# mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM22D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X881 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D12 io_analog[3] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X882 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X883 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X884 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X885 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X886 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X887 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X888 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X889 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X890 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X891 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X892 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X893 mpw5_submission_1/eigth_mirror_0/I_In mpw5_submission_1/isource_0/VM22D a_171016_648702# vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X894 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X895 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X896 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X897 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X898 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X899 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X900 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X901 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X902 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X903 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X904 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X905 mpw5_submission_0/eigth_mirror_0/I_out_4 mpw5_submission_0/eigth_mirror_0/I_In a_429020_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X906 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X907 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X908 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X909 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X910 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X911 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X912 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X913 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X914 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X915 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X916 a_433070_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X917 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X918 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X919 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X920 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X921 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X922 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X923 a_189936_651879# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X924 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X925 a_186120_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X926 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X927 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X928 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X929 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X930 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X931 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X932 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X933 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X934 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X935 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X936 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X937 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X938 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X939 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X940 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X941 a_430370_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X942 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X943 a_441658_643680# mpw5_submission_0/cmirror_channel_0/I_in_channel vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X944 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X945 mpw5_submission_1/tia_core_0/VM5D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 io_analog[6] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X946 mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X947 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X948 vssd1 mpw5_submission_1/cmirror_channel_0/I_in_channel sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X949 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X950 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X951 mpw5_submission_0/cmirror_channel_0/I_in_channel mpw5_submission_0/cmirror_channel_0/I_in_channel a_440818_643680# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X952 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X953 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X954 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X955 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X956 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X957 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X958 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X959 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X960 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X961 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X962 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X963 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X964 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X965 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X966 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X967 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X968 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X969 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X970 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X971 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X972 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X973 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X974 vccd1 mpw5_submission_1/outd_0/V_da2_N vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X975 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X976 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X977 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X978 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X979 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X980 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X981 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X982 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X983 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X984 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X985 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X986 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X987 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X988 a_443850_641883# a_441720_645346# mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X989 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X990 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X991 vccd1 io_analog[4] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X992 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X993 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X994 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X995 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X996 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X997 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X998 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X999 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1000 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1001 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1002 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1003 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1004 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1005 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1006 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_195570_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1007 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1008 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1009 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1010 mpw5_submission_1/tia_core_0/Out_2 mpw5_submission_1/outd_0/InputSignal io_analog[6] io_analog[6] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1011 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1012 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1013 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1014 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1015 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1016 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1017 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1018 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1019 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1020 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1021 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1022 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1023 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM6D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1024 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1025 mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__cap_var_lvt pd=0u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X1026 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1027 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1028 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1029 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1030 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1031 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1032 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1033 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1034 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1035 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1036 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1037 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1038 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1039 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1040 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1041 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1042 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1043 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1044 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1045 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1046 mpw5_submission_1/isource_0/VM22D a_171016_648702# mpw5_submission_1/isource_0/VM3D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1047 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1048 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1049 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1050 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1051 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1052 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1053 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1054 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1055 mpw5_submission_1/isource_0/VM12G mpw5_submission_1/isource_0/VM14D vccd1 mpw5_submission_1/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1056 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1057 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1058 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1059 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1060 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1061 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1062 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1063 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1064 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1065 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1066 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1067 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1068 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1069 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1070 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1071 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1072 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1073 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1074 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1075 a_464438_656600# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1076 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1077 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1078 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1079 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1080 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1081 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1082 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1083 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1084 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1085 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1086 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1087 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1088 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1089 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1090 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1091 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1092 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1093 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1094 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1095 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1096 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1097 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1098 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1099 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1100 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1101 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1102 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1103 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1104 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1105 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1106 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1107 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1108 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1109 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1110 a_431720_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1111 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1112 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1113 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1114 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1115 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1116 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1117 io_analog[3] mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/tia_core_0/Out_2 io_analog[3] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1118 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1119 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1120 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1121 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1122 vssd1 mpw5_submission_1/isource_0/VM12G mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1123 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1124 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1125 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1126 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1127 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1128 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1129 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1130 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1131 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1132 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1133 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1134 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1135 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1136 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1137 vccd1 mpw5_submission_0/isource_0/VM14D mpw5_submission_0/isource_0/VM12G mpw5_submission_0/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1138 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1139 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1140 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1141 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1142 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1143 a_201458_647480# mpw5_submission_1/cmirror_channel_0/I_in_channel vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1144 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1145 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1146 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1147 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1148 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1149 mpw5_submission_1/tia_core_0/VM31D mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1150 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1151 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1152 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1153 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1154 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1155 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1156 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1157 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1158 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1159 vccd1 mpw5_submission_1/isource_0/VM8D sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X1160 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1161 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1162 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1163 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1164 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1165 vccd1 io_analog[4] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1166 mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1167 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1168 mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1169 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1170 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1171 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1172 mpw5_submission_0/outd_0/V_da2_N vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1173 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1174 a_430370_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1175 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1176 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1177 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1178 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1179 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1180 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1181 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1182 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1183 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_657119# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1184 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1185 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1186 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1187 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1188 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1189 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1190 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1191 a_433070_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1192 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1193 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1194 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1195 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1196 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1197 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1198 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1199 a_186120_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1200 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1201 mpw5_submission_1/isource_0/VM3G a_185326_655038# vssd1 sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X1202 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1203 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1204 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1205 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1206 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1207 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1208 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1209 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1210 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1211 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1212 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1213 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1214 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
D13 vssd1 io_analog[7] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X1215 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1216 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1217 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1218 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1219 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1220 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1221 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1222 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1223 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1224 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1225 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1226 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1227 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1228 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1229 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1230 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D14 io_analog[2] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X1231 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1232 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1233 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1234 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D15 vssd1 io_analog[0] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X1235 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1236 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1237 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1238 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1239 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1240 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1241 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1242 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1243 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1244 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1245 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1246 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1247 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1248 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1249 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1250 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1251 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1252 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1253 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1254 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1255 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1256 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1257 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1258 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1259 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1260 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1261 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1262 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1263 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_429020_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1264 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1265 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1266 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1267 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1268 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1269 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1270 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1271 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1272 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1273 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1274 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1275 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1276 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1277 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1278 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1279 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1280 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1281 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1282 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1283 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1284 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1285 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM31D mpw5_submission_0/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1286 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1287 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1288 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1289 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1290 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1291 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1292 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1293 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1294 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1295 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1296 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1297 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1298 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1299 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1300 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1301 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1302 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1303 mpw5_submission_1/eigth_mirror_0/I_out_4 mpw5_submission_1/eigth_mirror_0/I_In a_188820_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1304 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1305 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1306 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1307 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1308 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1309 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1310 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_427670_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1311 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1312 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1313 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1314 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1315 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1316 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1317 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1318 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1319 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1320 a_430136_648079# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1321 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1322 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1323 vssd1 mpw5_submission_1/cmirror_channel_0/I_in_channel a_200618_647480# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1324 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1325 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1326 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1327 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1328 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1329 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1330 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1331 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1332 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1333 io_analog[1] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1334 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1335 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1336 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1337 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1338 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1339 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1340 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1341 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1342 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1343 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1344 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1345 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1346 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1347 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1348 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1349 mpw5_submission_0/isource_0/VM22D a_411216_644902# mpw5_submission_0/isource_0/VM3D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1350 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1351 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM12G vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1352 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1353 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1354 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1355 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1356 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1357 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1358 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1359 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1360 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1361 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1362 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1363 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_429020_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1364 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1365 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1366 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1367 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1368 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_426320_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1369 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/InputRef mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1370 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1371 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1372 a_429646_642496# a_430176_644928# vssd1 sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X1373 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1374 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1375 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1376 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1377 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1378 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1379 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1380 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1381 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1382 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1383 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1384 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1385 mpw5_submission_0/isource_0/VM12G mpw5_submission_0/isource_0/VM14D vccd1 mpw5_submission_0/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1386 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1387 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM31D mpw5_submission_1/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1388 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1389 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1390 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1391 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1392 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1393 mpw5_submission_1/tia_core_0/Out_2 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1394 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1395 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1396 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1397 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1398 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1399 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1400 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1401 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1402 mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/InputRef mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1403 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1404 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1405 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1406 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1407 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1408 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1409 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1410 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1411 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1412 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1413 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1414 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1415 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1416 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1417 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1418 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1419 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1420 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1421 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1422 mpw5_submission_0/tia_core_0/VM31D vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1423 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1424 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1425 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1426 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1427 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1428 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1429 a_201720_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1430 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1431 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1432 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1433 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1434 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1435 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1436 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1437 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1438 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1439 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1440 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1441 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1442 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1443 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1444 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1445 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1446 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1447 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1448 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1449 a_203370_649243# a_201520_649146# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1450 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1451 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1452 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1453 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1454 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1455 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1456 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1457 mpw5_submission_1/tia_core_0/VM31D mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1458 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1459 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1460 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1461 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1462 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1463 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1464 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1465 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1466 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1467 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1468 a_190170_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1469 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1470 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM31D mpw5_submission_1/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1471 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1472 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1473 mpw5_submission_0/tia_core_0/Out_2 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1474 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1475 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1476 mpw5_submission_0/outd_0/InputSignal io_analog[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1477 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1478 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1479 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1480 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1481 vssd1 vccd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1482 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1483 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1484 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1485 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1486 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1487 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1488 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1489 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1490 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1491 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1492 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1493 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1494 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1495 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1496 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1497 a_430370_636823# mpw5_submission_0/eigth_mirror_0/I_In mpw5_submission_0/eigth_mirror_0/I_out_3 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1498 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1499 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1500 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1501 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1502 mpw5_submission_0/tia_core_0/VM31D mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1503 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1504 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1505 vccd1 a_441720_645346# a_441920_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1506 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1507 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1508 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1509 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1510 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1511 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1512 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1513 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1514 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1515 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1516 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1517 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1518 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1519 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1520 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1521 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1522 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1523 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1524 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1525 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1526 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1527 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1528 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1529 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1530 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1531 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1532 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1533 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1534 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1535 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1536 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1537 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1538 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1539 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1540 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1541 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1542 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/InputRef mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1543 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1544 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1545 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1546 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1547 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1548 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1549 mpw5_submission_1/outd_0/V_da1_P vccd1 vssd1 sky130_fd_pr__res_high_po_2p85 l=6e+06u
X1550 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1551 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1552 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1553 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1554 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1555 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1556 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1557 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1558 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1559 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1560 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1561 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1562 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1563 a_426056_648806# a_426586_651238# vssd1 sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X1564 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1565 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1566 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1567 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1568 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM31D mpw5_submission_0/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1569 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1570 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1571 vssd1 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1572 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1573 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1574 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1575 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1576 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1577 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1578 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1579 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1580 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1581 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1582 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1583 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1584 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1585 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1586 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1587 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1588 a_429020_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1589 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1590 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1591 mpw5_submission_0/tia_core_0/VM31D mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1592 io_analog[0] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1593 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1594 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1595 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1596 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1597 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1598 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1599 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1600 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1601 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1602 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1603 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1604 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1605 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1606 a_443570_645443# a_441720_645346# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1607 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1608 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1609 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1610 mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1611 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1612 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1613 a_426320_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1614 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1615 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1616 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1617 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1618 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1619 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1620 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1621 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1622 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1623 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1624 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1625 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1626 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1627 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1628 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1629 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1630 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1631 vccd1 io_analog[1] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1632 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1633 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1634 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1635 a_189936_651879# mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM14D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X1636 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1637 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1638 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1639 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1640 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1641 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1642 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1643 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1644 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1645 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1646 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1647 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1648 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1649 a_171016_648702# mpw5_submission_1/isource_0/VM22D mpw5_submission_1/eigth_mirror_0/I_In vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1650 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1651 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1652 vccd1 io_analog[4] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1653 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1654 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1655 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1656 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1657 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1658 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1659 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1660 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1661 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1662 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1663 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_435770_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1664 a_443850_641883# a_441720_645346# mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1665 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1666 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1667 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1668 a_443570_645443# a_441720_645346# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1669 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1670 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1671 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1672 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1673 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1674 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1675 a_424970_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1676 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1677 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1678 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1679 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1680 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1681 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1682 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1683 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1684 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1685 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1686 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1687 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1688 a_189936_651879# mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM14D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X1689 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1690 a_189936_660919# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1691 a_203650_645683# a_201520_649146# mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1692 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1693 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1694 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1695 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1696 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1697 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1698 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1699 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1700 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1701 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1702 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1703 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1704 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1705 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1706 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1707 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1708 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1709 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM36D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1710 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1711 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1712 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1713 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1714 vssd1 mpw5_submission_1/cmirror_channel_0/I_in_channel a_202298_647480# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1715 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1716 a_201720_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1717 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1718 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1719 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1720 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1721 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1722 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1723 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1724 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1725 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1726 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1727 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1728 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1729 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1730 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1731 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1732 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1733 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1734 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1735 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1736 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1737 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1738 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1739 a_441920_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1740 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1741 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1742 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1743 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1744 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1745 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1746 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1747 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1748 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1749 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1750 a_430370_636823# mpw5_submission_0/eigth_mirror_0/I_In mpw5_submission_0/eigth_mirror_0/I_out_3 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1751 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1752 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1753 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1754 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1755 a_203370_649243# a_201520_649146# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1756 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1757 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1758 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1759 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1760 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1761 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1762 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1763 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1764 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1765 a_430136_654859# mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM8D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X1766 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1767 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1768 a_189936_651879# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1769 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1770 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1771 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1772 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1773 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1774 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1775 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1776 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1777 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1778 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1779 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1780 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1781 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1782 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1783 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1784 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1785 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_645809# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1786 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1787 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1788 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_657119# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1789 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1790 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1791 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1792 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1793 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1794 io_analog[6] mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/tia_core_0/Out_2 io_analog[6] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1795 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1796 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1797 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1798 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1799 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1800 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1801 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1802 mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1803 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1804 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1805 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1806 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1807 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1808 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1809 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1810 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1811 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1812 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1813 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1814 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1815 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1816 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1817 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1818 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1819 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1820 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1821 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1822 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1823 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1824 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1825 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1826 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1827 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1828 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1829 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1830 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1831 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_192870_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1832 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1833 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1834 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1835 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1836 a_171016_648702# mpw5_submission_1/isource_0/VM22D mpw5_submission_1/eigth_mirror_0/I_In vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1837 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1838 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1839 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1840 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1841 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1842 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1843 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1844 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1845 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1846 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1847 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1848 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1849 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1850 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1851 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1852 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1853 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1854 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1855 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1856 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1857 a_426320_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1858 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1859 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1860 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1861 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1862 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1863 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1864 a_430136_648079# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1865 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1866 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1867 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1868 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1869 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1870 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1871 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1872 a_429020_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1873 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1874 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1875 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1876 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1877 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1878 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1879 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1880 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1881 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_194220_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1882 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1883 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1884 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1885 mpw5_submission_0/tia_core_0/VM6D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1886 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1887 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1888 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1889 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1890 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1891 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1892 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1893 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1894 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1895 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1896 a_430370_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1897 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1898 mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1899 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1900 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1901 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1902 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1903 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1904 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1905 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1906 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1907 vccd1 io_analog[0] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1908 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1909 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1910 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1911 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1912 vssd1 vccd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1913 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1914 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1915 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1916 mpw5_submission_0/outd_0/V_da1_P vccd1 vssd1 sky130_fd_pr__res_high_po_2p85 l=6e+06u
X1917 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1918 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1919 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1920 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1921 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1922 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1923 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1924 a_427670_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1925 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1926 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1927 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1928 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1929 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1930 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1931 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1932 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1933 a_443570_645443# a_441720_645346# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1934 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1935 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1936 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1937 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1938 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1939 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1940 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1941 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1942 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1943 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1944 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1945 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1946 io_analog[0] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1947 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1948 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1949 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1950 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1951 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1952 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1953 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1954 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1955 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1956 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1957 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1958 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1959 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1960 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1961 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1962 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1963 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
D16 vssd1 io_analog[0] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X1964 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1965 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1966 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1967 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1968 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_658659# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1969 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1970 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1971 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_649609# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1972 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1973 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1974 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1975 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1976 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_195570_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1977 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1978 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1979 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1980 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1981 mpw5_submission_1/isource_0/VM22D a_171016_648702# mpw5_submission_1/isource_0/VM3D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1982 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1983 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1984 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1985 io_analog[1] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1986 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1987 mpw5_submission_0/isource_0/VM3D a_411216_644902# mpw5_submission_0/isource_0/VM22D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1988 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1989 a_189936_651879# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1990 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1991 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1992 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1993 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1994 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1995 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1996 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1997 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1998 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1999 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2000 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2001 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2002 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2003 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2004 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2005 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2006 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D17 io_analog[3] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X2007 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2008 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2009 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2010 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2011 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2012 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2013 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2014 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2015 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2016 mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2017 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2018 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2019 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2020 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2021 a_189936_649609# mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM22D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X2022 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2023 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2024 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2025 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2026 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2027 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2028 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2029 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2030 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2031 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2032 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2033 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2034 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2035 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2036 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2037 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2038 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2039 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2040 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2041 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2042 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2043 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2044 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2045 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2046 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2047 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2048 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2049 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2050 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2051 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2052 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2053 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2054 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2055 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2056 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2057 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2058 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2059 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2060 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2061 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2062 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2063 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2064 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2065 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2066 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2067 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2068 mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2069 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2070 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2071 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2072 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2073 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2074 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2075 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2076 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_192870_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2077 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2078 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2079 mpw5_submission_0/tia_core_0/VM6D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2080 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2081 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2082 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X2083 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2084 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2085 vssd1 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM36D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2086 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2087 a_184770_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2088 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2089 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2090 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2091 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2092 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2093 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2094 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2095 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2096 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2097 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2098 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2099 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2100 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2101 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2102 vccd1 mpw5_submission_0/outd_0/V_da2_P vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2103 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2104 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_190170_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2105 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2106 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2107 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2108 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2109 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2110 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2111 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2112 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2113 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2114 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2115 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2116 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2117 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2118 mpw5_submission_1/tia_core_0/Out_2 mpw5_submission_1/outd_0/InputSignal io_analog[6] io_analog[6] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2119 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2120 mpw5_submission_0/isource_0/VM22D a_411216_644902# mpw5_submission_0/isource_0/VM3D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X2121 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2122 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2123 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2124 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2125 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2126 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2127 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2128 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2129 mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2130 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2131 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2132 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2133 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2134 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2135 mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/InputRef mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2136 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2137 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2138 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2139 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2140 io_analog[0] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2141 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2142 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2143 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2144 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2145 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2146 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2147 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2148 a_195570_640623# mpw5_submission_1/eigth_mirror_0/I_In mpw5_submission_1/eigth_mirror_0/I_In vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2149 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2150 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2151 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2152 vccd1 mpw5_submission_0/isource_0/VM14D mpw5_submission_0/isource_0/VM12G mpw5_submission_0/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2153 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2154 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2155 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2156 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2157 mpw5_submission_1/outd_0/InputSignal io_analog[6] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2158 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2159 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2160 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2161 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2162 a_433070_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2163 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2164 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2165 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2166 vssd1 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X2167 io_analog[1] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2168 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2169 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2170 vssd1 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X2171 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2172 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2173 a_186120_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2174 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2175 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2176 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2177 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2178 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2179 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2180 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2181 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2182 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2183 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2184 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2185 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2186 a_443570_645443# a_441720_645346# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2187 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2188 mpw5_submission_1/tia_core_0/VM36D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM39D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2189 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2190 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2191 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2192 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2193 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2194 mpw5_submission_1/isource_0/VM3D a_171016_648702# mpw5_submission_1/isource_0/VM22D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X2195 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2196 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2197 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2198 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2199 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2200 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2201 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2202 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2203 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X2204 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2205 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2206 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2207 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2208 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2209 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2210 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2211 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2212 a_194220_640623# mpw5_submission_1/eigth_mirror_0/I_In mpw5_submission_1/cmirror_channel_0/I_in_channel vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2213 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2214 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2215 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2216 a_431720_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2217 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2218 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2219 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2220 a_440818_643680# mpw5_submission_0/cmirror_channel_0/I_in_channel vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2221 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2222 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2223 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2224 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2225 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2226 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2227 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2228 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2229 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2230 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2231 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2232 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2233 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2234 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2235 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2236 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2237 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2238 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2239 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2240 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2241 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2242 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2243 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2244 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2245 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2246 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2247 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2248 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2249 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2250 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2251 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2252 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2253 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM31D mpw5_submission_1/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2254 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2255 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2256 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2257 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2258 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2259 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2260 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2261 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2262 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2263 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2264 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2265 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2266 a_430370_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2267 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2268 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2269 vccd1 a_201520_649146# a_201720_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2270 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2271 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2272 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2273 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2274 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2275 vccd1 vssd1 mpw5_submission_1/tia_core_0/VM31D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2276 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2277 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2278 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2279 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2280 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2281 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2282 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2283 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2284 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2285 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2286 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2287 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2288 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2289 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2290 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2291 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2292 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2293 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2294 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2295 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2296 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2297 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2298 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2299 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2300 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2301 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2302 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2303 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2304 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D18 io_analog[7] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X2305 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2306 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2307 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2308 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2309 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2310 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2311 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2312 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2313 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2314 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2315 a_189936_651879# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2316 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2317 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2318 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2319 vssd1 mpw5_submission_0/isource_0/VM3G mpw5_submission_0/isource_0/VM3D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X2320 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2321 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2322 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2323 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2324 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2325 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2326 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2327 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2328 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2329 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2330 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2331 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2332 a_443850_641883# a_441720_645346# mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2333 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2334 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2335 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2336 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2337 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2338 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2339 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2340 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2341 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2342 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2343 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2344 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2345 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2346 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2347 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2348 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2349 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2350 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2351 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2352 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2353 a_443570_645443# a_441720_645346# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2354 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2355 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2356 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM6D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2357 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2358 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2359 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2360 a_441658_643680# mpw5_submission_0/cmirror_channel_0/I_in_channel vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2361 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2362 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2363 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2364 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2365 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2366 mpw5_submission_0/tia_core_0/VM31D mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2367 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2368 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2369 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2370 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2371 a_430136_648079# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2372 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2373 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D19 io_analog[3] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X2374 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2375 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2376 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2377 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2378 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2379 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2380 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2381 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2382 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2383 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2384 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2385 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2386 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2387 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2388 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2389 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2390 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2391 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2392 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2393 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_645809# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2394 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2395 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2396 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2397 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2398 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2399 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2400 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2401 mpw5_submission_1/eigth_mirror_0/I_out_4 mpw5_submission_1/eigth_mirror_0/I_In a_188820_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2402 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2403 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2404 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2405 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2406 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2407 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2408 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2409 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2410 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2411 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2412 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2413 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2414 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2415 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2416 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2417 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2418 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2419 mpw5_submission_1/eigth_mirror_0/I_In mpw5_submission_1/isource_0/VM22D a_171016_648702# vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2420 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2421 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2422 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2423 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2424 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2425 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2426 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2427 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2428 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2429 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2430 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2431 mpw5_submission_0/outd_0/InputSignal io_analog[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2432 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2433 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2434 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2435 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2436 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2437 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2438 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2439 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2440 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2441 mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2442 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2443 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2444 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2445 io_analog[0] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2446 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2447 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2448 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2449 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2450 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2451 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2452 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2453 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2454 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2455 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2456 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2457 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2458 vccd1 a_201520_649146# a_201720_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2459 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2460 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2461 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2462 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2463 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2464 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2465 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2466 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2467 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2468 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2469 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2470 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2471 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2472 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2473 vccd1 io_analog[1] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2474 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2475 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2476 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2477 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2478 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2479 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2480 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2481 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2482 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2483 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2484 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2485 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2486 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2487 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2488 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2489 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2490 a_424970_636823# mpw5_submission_0/eigth_mirror_0/I_In mpw5_submission_0/eigth_mirror_0/I_out_7 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2491 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2492 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2493 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2494 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2495 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2496 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2497 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2498 vssd1 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 sky130_fd_pr__cap_mim_m3_1 l=1.2e+07u w=1.5e+07u
X2499 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2500 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2501 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2502 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2503 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2504 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2505 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2506 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2507 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2508 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2509 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2510 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2511 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2512 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2513 vssd1 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X2514 a_189446_646296# a_189976_648728# vssd1 sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X2515 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2516 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2517 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2518 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2519 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2520 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2521 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2522 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2523 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2524 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2525 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2526 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2527 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2528 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2529 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2530 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2531 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2532 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2533 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2534 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2535 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2536 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2537 mpw5_submission_0/isource_0/VM3D mpw5_submission_0/isource_0/VM3G vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X2538 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2539 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2540 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2541 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2542 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2543 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2544 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2545 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2546 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D20 vssd1 io_analog[0] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X2547 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2548 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2549 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2550 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2551 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2552 mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2553 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2554 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2555 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2556 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2557 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D21 vssd1 io_analog[2] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
D22 vssd1 io_analog[1] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X2558 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2559 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2560 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2561 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2562 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2563 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2564 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2565 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2566 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2567 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2568 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2569 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2570 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2571 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2572 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2573 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2574 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2575 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2576 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2577 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2578 mpw5_submission_1/tia_core_0/VM31D mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2579 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2580 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2581 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2582 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2583 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2584 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2585 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2586 a_187470_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2587 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2588 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2589 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2590 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2591 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2592 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2593 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2594 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2595 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2596 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2597 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2598 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2599 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X2600 a_426320_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2601 mpw5_submission_0/outd_0/InputSignal io_analog[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2602 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2603 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2604 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2605 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2606 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2607 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2608 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2609 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2610 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2611 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2612 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2613 mpw5_submission_1/eigth_mirror_0/I_In mpw5_submission_1/isource_0/VM22D a_171016_648702# vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2614 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2615 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2616 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2617 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_195570_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2618 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2619 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2620 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2621 mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/InputRef mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2622 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2623 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2624 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2625 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2626 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2627 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2628 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2629 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2630 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2631 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2632 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2633 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2634 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2635 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2636 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2637 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2638 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2639 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2640 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2641 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2642 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2643 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2644 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2645 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2646 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2647 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2648 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_188820_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2649 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2650 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2651 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2652 io_analog[5] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2653 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2654 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2655 vccd1 mpw5_submission_1/isource_0/VM14D mpw5_submission_1/isource_0/VM12G mpw5_submission_1/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2656 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2657 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2658 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2659 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2660 a_424970_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2661 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2662 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2663 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2664 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2665 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2666 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2667 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2668 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2669 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2670 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2671 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2672 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2673 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2674 vccd1 mpw5_submission_0/outd_0/V_da2_N vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2675 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2676 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2677 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2678 mpw5_submission_0/tia_core_0/VM36D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM39D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2679 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_194220_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2680 mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2681 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2682 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2683 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2684 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2685 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2686 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2687 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2688 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2689 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2690 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2691 vssd1 vccd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2692 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_654859# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2693 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2694 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2695 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2696 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2697 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2698 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2699 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2700 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2701 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2702 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM31D mpw5_submission_0/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2703 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2704 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2705 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2706 mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2707 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2708 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2709 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2710 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2711 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2712 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2713 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2714 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2715 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2716 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2717 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2718 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2719 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2720 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2721 mpw5_submission_1/eigth_mirror_0/I_In mpw5_submission_1/isource_0/VM22D a_171016_648702# vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2722 mpw5_submission_1/tia_core_0/VM6D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2723 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2724 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2725 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2726 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2727 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2728 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2729 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2730 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X2731 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2732 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2733 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D23 vssd1 io_analog[3] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X2734 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2735 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2736 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2737 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2738 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2739 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2740 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2741 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2742 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2743 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X2744 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2745 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2746 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2747 vccd1 vssd1 mpw5_submission_0/tia_core_0/Out_2 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2748 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2749 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2750 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X2751 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2752 vccd1 vssd1 mpw5_submission_1/tia_core_0/Out_2 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2753 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2754 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2755 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2756 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2757 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2758 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2759 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2760 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2761 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2762 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2763 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2764 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2765 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2766 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2767 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2768 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2769 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2770 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2771 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2772 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_435770_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2773 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2774 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2775 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2776 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2777 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2778 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2779 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2780 a_442498_643680# mpw5_submission_0/cmirror_channel_0/I_in_channel mpw5_submission_0/cmirror_channel_0/TIA_I_Bias2 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2781 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_430370_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2782 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2783 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2784 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2785 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2786 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2787 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2788 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2789 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2790 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2791 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2792 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_433070_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2793 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2794 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2795 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2796 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_430370_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2797 vssd1 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 sky130_fd_pr__cap_mim_m3_1 l=1.2e+07u w=1.5e+07u
X2798 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2799 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2800 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2801 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2802 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2803 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2804 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2805 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2806 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2807 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2808 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2809 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2810 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2811 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2812 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2813 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2814 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2815 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2816 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2817 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2818 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2819 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2820 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2821 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2822 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2823 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2824 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2825 a_189936_651879# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2826 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2827 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2828 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2829 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2830 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2831 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2832 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2833 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2834 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2835 io_analog[5] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2836 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2837 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2838 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2839 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2840 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2841 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2842 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2843 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2844 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2845 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2846 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2847 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2848 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_431720_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2849 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2850 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2851 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2852 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_184770_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2853 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2854 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2855 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2856 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2857 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM6D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2858 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2859 a_429020_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2860 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2861 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2862 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2863 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2864 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2865 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2866 mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2867 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2868 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2869 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2870 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2871 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2872 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2873 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2874 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2875 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2876 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2877 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2878 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2879 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2880 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2881 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2882 vssd1 mpw5_submission_0/isource_0/VM11D a_422158_661070# vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X2883 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2884 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2885 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2886 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2887 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2888 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2889 mpw5_submission_1/isource_0/VM12G mpw5_submission_1/isource_0/VM14D vccd1 mpw5_submission_1/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2890 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2891 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2892 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2893 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2894 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2895 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2896 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2897 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2898 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2899 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2900 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2901 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2902 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2903 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2904 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2905 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2906 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2907 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2908 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2909 a_427670_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2910 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2911 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2912 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2913 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2914 a_189936_658659# mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM8D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X2915 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2916 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2917 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2918 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2919 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2920 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D24 vssd1 io_analog[2] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X2921 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2922 a_430136_648079# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2923 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2924 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2925 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2926 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2927 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2928 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2929 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2930 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2931 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2932 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2933 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2934 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2935 mpw5_submission_0/outd_0/V_da1_N vccd1 vssd1 sky130_fd_pr__res_high_po_2p85 l=6e+06u
X2936 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2937 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2938 a_428176_648806# a_428706_651238# vssd1 sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X2939 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2940 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2941 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2942 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2943 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2944 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X2945 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2946 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2947 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM36D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2948 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2949 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2950 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2951 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2952 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2953 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2954 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2955 a_426320_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2956 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2957 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2958 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2959 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2960 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2961 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2962 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2963 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2964 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2965 mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2966 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2967 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2968 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2969 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2970 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2971 mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2972 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2973 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2974 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2975 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X2976 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2977 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2978 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2979 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2980 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2981 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2982 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2983 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2984 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D25 io_analog[3] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X2985 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2986 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2987 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2988 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2989 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2990 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2991 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2992 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2993 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2994 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2995 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2996 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2997 a_190170_640623# mpw5_submission_1/eigth_mirror_0/I_In mpw5_submission_1/eigth_mirror_0/I_out_3 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2998 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2999 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3000 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3001 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3002 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3003 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3004 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3005 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3006 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3007 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3008 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3009 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3010 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3011 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3012 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3013 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3014 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3015 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3016 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3017 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D26 vssd1 io_analog[2] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X3018 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3019 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3020 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3021 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3022 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3023 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3024 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3025 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3026 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3027 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3028 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3029 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3030 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3031 vssd1 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM6D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3032 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3033 a_443570_645443# a_441720_645346# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3034 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3035 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3036 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3037 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3038 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3039 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3040 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3041 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3042 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3043 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3044 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3045 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3046 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3047 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3048 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3049 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3050 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3051 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3052 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3053 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3054 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3055 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3056 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3057 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X3058 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM36D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3059 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3060 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3061 a_203650_645683# a_201520_649146# mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3062 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3063 vssd1 mpw5_submission_1/isource_0/VM3G mpw5_submission_1/isource_0/VM3D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3064 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3065 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3066 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3067 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3068 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3069 a_430136_648079# mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM14D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X3070 mpw5_submission_1/isource_0/VM12G mpw5_submission_1/isource_0/VM14D vccd1 mpw5_submission_1/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3071 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3072 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3073 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3074 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3075 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_190170_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3076 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3077 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3078 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3079 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3080 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3081 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3082 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3083 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3084 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3085 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3086 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3087 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/InputRef mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3088 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3089 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3090 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3091 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3092 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3093 a_443850_641883# a_441720_645346# mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3094 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3095 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3096 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3097 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
D27 vssd1 io_analog[8] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X3098 a_441920_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3099 mpw5_submission_1/outd_0/InputSignal io_analog[6] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3100 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3101 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3102 mpw5_submission_0/isource_0/VM12G mpw5_submission_0/isource_0/VM14D vccd1 mpw5_submission_0/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3103 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3104 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3105 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3106 io_analog[4] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3107 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3108 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3109 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3110 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3111 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3112 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3113 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3114 a_203650_645683# a_201520_649146# mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3115 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3116 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3117 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3118 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3119 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3120 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D28 io_analog[1] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X3121 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3122 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3123 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3124 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3125 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3126 mpw5_submission_1/tia_core_0/VM6D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3127 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3128 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3129 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3130 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3131 vccd1 io_analog[5] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3132 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3133 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3134 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3135 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3136 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3137 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3138 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3139 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3140 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3141 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3142 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3143 mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3144 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3145 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3146 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3147 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3148 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3149 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3150 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3151 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3152 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3153 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3154 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D29 vssd1 io_analog[7] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X3155 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3156 a_431720_636823# mpw5_submission_0/eigth_mirror_0/I_In mpw5_submission_0/eigth_mirror_0/I_out_2 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3157 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3158 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3159 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3160 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3161 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3162 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3163 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3164 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3165 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3166 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3167 mpw5_submission_1/outd_0/V_da2_P vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3168 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3169 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3170 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3171 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3172 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3173 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3174 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3175 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3176 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3177 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3178 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3179 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3180 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3181 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3182 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3183 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3184 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3185 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3186 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3187 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3188 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3189 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3190 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3191 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3192 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3193 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3194 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3195 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3196 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3197 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3198 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3199 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3200 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3201 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3202 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3203 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3204 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3205 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3206 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3207 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3208 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3209 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3210 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3211 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3212 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3213 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3214 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3215 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3216 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3217 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3218 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3219 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3220 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3221 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3222 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3223 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3224 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3225 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3226 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM36D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3227 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3228 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3229 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3230 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3231 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3232 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3233 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3234 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3235 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3236 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3237 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3238 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3239 vccd1 io_analog[5] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3240 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3241 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3242 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3243 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3244 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3245 mpw5_submission_1/outd_0/InputSignal io_analog[6] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3246 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3247 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3248 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3249 mpw5_submission_1/isource_0/VM22D a_171016_648702# mpw5_submission_1/isource_0/VM3D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3250 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3251 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3252 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3253 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3254 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3255 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3256 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3257 mpw5_submission_1/isource_0/VM3D mpw5_submission_1/isource_0/VM3G vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3258 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3259 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3260 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3261 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3262 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_435770_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3263 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3264 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3265 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3266 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3267 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3268 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3269 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3270 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_660919# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3271 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_649609# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3272 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3273 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3274 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3275 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3276 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3277 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3278 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3279 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3280 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3281 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3282 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3283 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3284 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3285 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3286 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3287 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3288 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3289 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3290 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3291 a_189936_660919# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3292 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3293 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3294 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3295 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3296 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3297 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3298 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3299 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3300 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3301 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3302 mpw5_submission_0/tia_core_0/VM5D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 io_analog[3] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3303 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3304 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3305 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3306 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3307 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3308 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3309 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3310 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3311 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3312 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3313 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3314 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_434420_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3315 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3316 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3317 mpw5_submission_1/outd_0/V_da1_P vccd1 vssd1 sky130_fd_pr__res_high_po_2p85 l=6e+06u
X3318 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3319 mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3320 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3321 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3322 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3323 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3324 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3325 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3326 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3327 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3328 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3329 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3330 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3331 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3332 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3333 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3334 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3335 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3336 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3337 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3338 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3339 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3340 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3341 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3342 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3343 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3344 a_203650_645683# a_201520_649146# mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3345 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3346 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM31D mpw5_submission_1/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3347 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3348 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3349 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3350 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3351 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3352 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3353 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3354 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3355 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3356 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3357 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3358 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3359 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3360 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3361 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3362 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3363 a_189936_651879# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3364 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3365 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3366 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3367 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3368 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3369 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3370 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3371 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3372 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3373 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3374 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3375 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3376 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3377 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3378 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3379 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3380 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3381 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3382 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3383 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3384 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3385 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3386 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3387 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3388 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3389 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3390 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3391 mpw5_submission_0/eigth_mirror_0/I_out_3 mpw5_submission_0/eigth_mirror_0/I_In a_430370_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3392 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3393 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3394 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3395 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3396 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3397 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3398 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3399 mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3400 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3401 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3402 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3403 vccd1 io_analog[4] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3404 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3405 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3406 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3407 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3408 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3409 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3410 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3411 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3412 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3413 mpw5_submission_1/tia_core_0/VM6D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3414 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3415 vccd1 io_analog[0] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3416 vssd1 vccd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3417 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM36D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3418 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3419 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3420 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3421 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3422 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3423 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3424 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3425 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3426 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3427 mpw5_submission_0/outd_0/InputSignal io_analog[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3428 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3429 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3430 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3431 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3432 io_analog[4] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3433 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3434 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3435 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3436 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3437 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3438 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3439 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3440 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3441 mpw5_submission_1/outd_0/V_da1_P vccd1 vssd1 sky130_fd_pr__res_high_po_2p85 l=6e+06u
X3442 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3443 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3444 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3445 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3446 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3447 vssd1 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3448 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3449 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3450 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3451 mpw5_submission_0/outd_0/InputSignal io_analog[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3452 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3453 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3454 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3455 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3456 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3457 io_analog[1] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3458 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3459 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3460 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3461 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3462 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3463 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3464 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3465 io_analog[5] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3466 mpw5_submission_1/isource_0/VM3D a_171016_648702# mpw5_submission_1/isource_0/VM22D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3467 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3468 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3469 a_191520_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3470 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3471 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3472 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3473 a_171016_648702# mpw5_submission_1/isource_0/VM22D mpw5_submission_1/eigth_mirror_0/I_In vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3474 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3475 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3476 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3477 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3478 vccd1 mpw5_submission_1/outd_0/V_da2_P vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3479 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3480 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3481 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3482 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3483 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3484 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3485 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3486 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3487 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3488 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3489 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D30 io_analog[2] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X3490 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3491 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3492 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3493 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3494 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3495 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3496 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3497 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3498 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3499 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3500 mpw5_submission_0/tia_core_0/Out_2 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3501 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3502 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3503 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3504 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D31 io_analog[3] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X3505 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3506 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3507 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3508 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3509 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3510 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3511 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3512 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3513 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3514 mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3515 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3516 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3517 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3518 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3519 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3520 mpw5_submission_1/tia_core_0/VM31D vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3521 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3522 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3523 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3524 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3525 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_427670_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3526 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3527 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3528 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3529 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3530 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3531 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3532 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3533 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3534 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3535 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3536 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3537 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3538 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3539 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3540 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3541 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3542 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3543 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3544 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3545 mpw5_submission_0/outd_0/InputSignal io_analog[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3546 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3547 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3548 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3549 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3550 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3551 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3552 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3553 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3554 mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3555 mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3556 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3557 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3558 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3559 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3560 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3561 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3562 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3563 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3564 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3565 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3566 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3567 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3568 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3569 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3570 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3571 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3572 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3573 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3574 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3575 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3576 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3577 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3578 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_195570_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3579 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3580 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3581 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3582 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3583 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3584 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3585 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3586 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3587 mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/InputRef mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3588 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3589 vssd1 a_428706_651238# vssd1 sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X3590 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3591 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3592 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3593 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3594 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3595 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3596 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3597 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3598 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3599 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3600 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3601 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3602 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3603 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3604 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3605 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3606 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3607 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3608 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3609 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3610 mpw5_submission_0/tia_core_0/VM31D vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3611 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3612 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3613 mpw5_submission_0/tia_core_0/VM6D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3614 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3615 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3616 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3617 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3618 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3619 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3620 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3621 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3622 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3623 mpw5_submission_0/isource_0/VM3D a_411216_644902# mpw5_submission_0/isource_0/VM22D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3624 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3625 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3626 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3627 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3628 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3629 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3630 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3631 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3632 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3633 a_186916_652606# a_186386_655038# vssd1 sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X3634 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3635 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_194220_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3636 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3637 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3638 io_analog[4] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3639 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3640 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3641 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3642 mpw5_submission_1/outd_0/InputSignal io_analog[6] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3643 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3644 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3645 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3646 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3647 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3648 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3649 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3650 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3651 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3652 vccd1 mpw5_submission_1/isource_0/VM14D mpw5_submission_1/isource_0/VM12G mpw5_submission_1/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3653 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3654 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3655 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3656 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3657 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3658 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3659 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3660 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3661 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3662 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3663 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3664 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3665 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3666 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3667 io_analog[5] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3668 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3669 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3670 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3671 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3672 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3673 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3674 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3675 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3676 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3677 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3678 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3679 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3680 mpw5_submission_1/tia_core_0/VM31D mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3681 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3682 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3683 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_192870_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3684 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3685 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3686 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3687 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3688 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3689 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3690 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3691 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3692 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3693 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3694 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3695 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3696 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3697 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3698 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3699 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3700 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3701 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3702 mpw5_submission_0/outd_0/V_da2_P vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3703 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3704 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3705 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3706 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3707 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3708 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3709 mpw5_submission_0/isource_0/VM8D a_422158_661070# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X3710 mpw5_submission_0/isource_0/VM3G a_424386_651238# vssd1 sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X3711 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3712 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3713 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3714 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3715 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3716 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3717 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3718 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3719 a_203370_649243# a_201520_649146# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3720 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3721 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3722 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3723 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3724 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3725 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3726 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3727 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3728 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3729 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3730 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3731 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3732 a_443570_645443# a_441720_645346# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3733 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3734 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3735 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3736 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3737 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3738 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3739 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3740 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3741 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3742 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3743 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3744 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3745 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3746 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3747 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3748 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_194220_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3749 mpw5_submission_1/outd_0/V_da2_N vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3750 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3751 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3752 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3753 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3754 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D32 vssd1 io_analog[1] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X3755 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3756 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3757 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3758 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3759 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3760 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3761 a_189936_651879# mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM14D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X3762 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3763 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_433070_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3764 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3765 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_430370_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3766 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3767 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias2 mpw5_submission_1/cmirror_channel_0/I_in_channel a_202298_647480# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3768 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3769 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3770 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3771 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3772 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3773 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3774 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3775 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3776 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3777 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3778 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3779 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3780 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3781 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3782 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3783 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3784 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3785 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3786 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3787 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3788 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3789 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3790 a_430136_654859# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3791 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3792 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3793 mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/InputRef mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3794 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3795 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3796 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3797 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3798 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3799 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3800 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3801 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3802 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3803 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3804 mpw5_submission_0/tia_core_0/VM36D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3805 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3806 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3807 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3808 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3809 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3810 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3811 a_195570_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3812 mpw5_submission_1/eigth_mirror_0/I_out_3 mpw5_submission_1/eigth_mirror_0/I_In a_190170_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3813 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3814 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3815 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3816 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3817 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3818 vssd1 a_431236_644928# vssd1 sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X3819 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3820 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3821 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3822 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3823 vssd1 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3824 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3825 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3826 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_431720_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3827 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3828 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3829 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3830 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D33 io_analog[7] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X3831 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3832 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3833 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3834 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3835 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_184770_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3836 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3837 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3838 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3839 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3840 mpw5_submission_0/outd_0/V_da1_P vccd1 vssd1 sky130_fd_pr__res_high_po_2p85 l=6e+06u
X3841 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3842 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3843 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3844 mpw5_submission_0/isource_0/VM3D mpw5_submission_0/isource_0/VM3G vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3845 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3846 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3847 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3848 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3849 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3850 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3851 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3852 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3853 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3854 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3855 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3856 vccd1 mpw5_submission_1/isource_0/VM14D mpw5_submission_1/isource_0/VM12G mpw5_submission_1/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3857 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3858 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3859 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3860 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3861 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3862 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3863 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3864 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3865 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3866 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3867 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3868 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3869 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3870 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3871 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3872 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3873 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3874 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3875 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3876 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3877 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3878 a_427670_636823# mpw5_submission_0/eigth_mirror_0/I_In mpw5_submission_0/eigth_mirror_0/I_out_5 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3879 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3880 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3881 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3882 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3883 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_430370_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3884 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3885 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3886 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3887 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3888 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3889 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3890 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3891 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3892 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3893 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3894 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3895 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3896 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3897 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3898 vccd1 a_201520_649146# a_201720_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3899 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3900 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3901 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3902 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3903 a_189936_651879# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3904 vccd1 mpw5_submission_0/outd_0/V_da2_N vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3905 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3906 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3907 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3908 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3909 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3910 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3911 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3912 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3913 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3914 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3915 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3916 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3917 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3918 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3919 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3920 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3921 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3922 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3923 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3924 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3925 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3926 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3927 a_426320_636823# mpw5_submission_0/eigth_mirror_0/I_In mpw5_submission_0/eigth_mirror_0/I_out_6 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3928 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3929 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3930 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3931 vssd1 mpw5_submission_1/cmirror_channel_0/I_in_channel a_202298_647480# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3932 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3933 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3934 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3935 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3936 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3937 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3938 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3939 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3940 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3941 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3942 mpw5_submission_0/outd_0/InputSignal io_analog[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3943 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3944 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3945 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3946 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3947 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3948 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3949 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3950 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3951 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3952 a_184770_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3953 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3954 vccd1 io_analog[5] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3955 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3956 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3957 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3958 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3959 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3960 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3961 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3962 io_analog[4] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3963 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3964 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3965 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3966 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3967 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3968 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3969 mpw5_submission_0/eigth_mirror_0/I_out_2 mpw5_submission_0/eigth_mirror_0/I_In a_431720_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3970 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3971 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3972 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3973 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3974 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3975 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3976 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3977 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3978 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3979 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3980 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3981 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3982 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3983 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3984 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3985 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3986 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3987 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3988 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3989 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3990 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3991 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3992 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3993 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3994 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3995 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
R0 vccd1 io_clamp_high[2] sky130_fd_pr__res_generic_m3 w=1.1e+07u l=250000u
X3996 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3997 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3998 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3999 a_430136_648079# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4000 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4001 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4002 a_184770_640623# mpw5_submission_1/eigth_mirror_0/I_In mpw5_submission_1/eigth_mirror_0/I_out_7 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4003 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4004 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4005 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4006 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4007 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4008 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4009 a_191520_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4010 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4011 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4012 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4013 io_analog[3] mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/tia_core_0/Out_2 io_analog[3] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4014 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4015 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4016 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4017 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4018 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4019 mpw5_submission_1/tia_core_0/VM36D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM39D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4020 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4021 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4022 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4023 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4024 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4025 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4026 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4027 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4028 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4029 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4030 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4031 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4032 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4033 a_443570_645443# a_441720_645346# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4034 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4035 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4036 vssd1 mpw5_submission_0/cmirror_channel_0/I_in_channel a_442498_643680# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4037 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4038 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4039 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4040 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4041 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4042 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4043 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4044 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4045 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4046 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4047 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4048 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4049 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4050 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4051 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4052 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4053 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4054 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4055 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4056 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4057 mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4058 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4059 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4060 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4061 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4062 a_201720_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4063 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4064 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4065 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4066 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4067 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4068 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4069 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4070 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4071 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4072 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4073 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4074 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4075 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4076 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4077 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4078 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4079 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4080 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4081 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4082 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4083 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4084 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4085 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4086 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4087 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4088 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4089 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4090 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4091 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4092 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4093 io_analog[3] mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM5D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4094 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4095 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4096 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4097 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4098 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4099 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4100 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4101 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4102 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4103 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4104 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4105 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4106 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4107 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4108 mpw5_submission_1/isource_0/VM22D a_171016_648702# mpw5_submission_1/isource_0/VM3D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4109 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4110 a_203650_645683# a_201520_649146# mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4111 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4112 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4113 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4114 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4115 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4116 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4117 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4118 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4119 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4120 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4121 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4122 vssd1 vccd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4123 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4124 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4125 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4126 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4127 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4128 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4129 a_430136_648079# mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM14D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X4130 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4131 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4132 mpw5_submission_1/outd_0/InputSignal io_analog[6] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4133 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4134 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4135 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4136 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4137 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4138 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4139 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4140 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4141 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4142 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4143 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4144 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4145 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4146 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4147 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4148 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4149 mpw5_submission_0/tia_core_0/VM5D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4150 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4151 io_analog[1] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4152 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4153 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4154 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4155 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4156 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4157 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4158 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4159 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_660919# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4160 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4161 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4162 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4163 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4164 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4165 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4166 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4167 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4168 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4169 vccd1 mpw5_submission_1/outd_0/V_da2_P vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4170 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4171 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4172 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4173 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4174 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4175 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4176 mpw5_submission_1/outd_0/V_da1_N vccd1 vssd1 sky130_fd_pr__res_high_po_2p85 l=6e+06u
X4177 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4178 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4179 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4180 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4181 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4182 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4183 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4184 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4185 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4186 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4187 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_658659# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4188 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4189 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4190 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4191 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4192 a_443850_641883# a_441720_645346# mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4193 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4194 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4195 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4196 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM6D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4197 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4198 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4199 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4200 io_analog[3] mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM5D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4201 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4202 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4203 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM6D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4204 mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4205 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4206 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4207 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4208 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4209 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4210 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4211 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4212 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4213 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4214 mpw5_submission_1/outd_0/InputSignal io_analog[6] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4215 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4216 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4217 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4218 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4219 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4220 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4221 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4222 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4223 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4224 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4225 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4226 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4227 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4228 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4229 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4230 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4231 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4232 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4233 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4234 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4235 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4236 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4237 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4238 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4239 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4240 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4241 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4242 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4243 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4244 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4245 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4246 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4247 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_188820_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4248 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4249 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4250 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4251 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4252 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4253 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4254 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4255 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4256 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4257 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4258 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4259 a_194220_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4260 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4261 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4262 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4263 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4264 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4265 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4266 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4267 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4268 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4269 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4270 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4271 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4272 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4273 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4274 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4275 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4276 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4277 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4278 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4279 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4280 mpw5_submission_1/tia_core_0/VM5D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 io_analog[6] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4281 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4282 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4283 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4284 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4285 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4286 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4287 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4288 a_186916_652606# a_187446_655038# vssd1 sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X4289 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4290 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4291 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4292 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4293 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4294 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4295 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4296 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4297 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4298 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4299 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4300 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4301 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D34 vssd1 io_analog[8] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X4302 mpw5_submission_1/outd_0/V_da1_N vccd1 vssd1 sky130_fd_pr__res_high_po_2p85 l=6e+06u
X4303 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4304 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4305 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4306 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4307 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4308 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4309 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4310 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4311 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4312 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4313 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4314 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4315 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4316 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4317 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4318 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4319 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4320 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4321 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4322 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4323 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4324 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4325 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4326 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4327 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4328 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4329 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4330 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4331 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4332 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4333 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4334 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4335 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4336 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4337 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4338 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4339 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4340 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4341 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4342 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4343 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4344 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4345 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4346 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4347 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4348 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4349 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4350 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4351 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4352 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4353 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4354 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4355 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4356 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4357 vssd1 mpw5_submission_1/isource_0/VM3G mpw5_submission_1/isource_0/VM3D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4358 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4359 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4360 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4361 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/InputRef mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4362 vccd1 vssd1 mpw5_submission_1/tia_core_0/Out_2 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D35 io_analog[2] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X4363 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4364 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4365 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4366 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_435770_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4367 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4368 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4369 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4370 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4371 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4372 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4373 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4374 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4375 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4376 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4377 mpw5_submission_0/outd_0/V_da2_P vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4378 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4379 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4380 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4381 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4382 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4383 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4384 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4385 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4386 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4387 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4388 mpw5_submission_0/outd_0/InputSignal io_analog[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4389 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4390 vssd1 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4391 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4392 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4393 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4394 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4395 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4396 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4397 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4398 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4399 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4400 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4401 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4402 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4403 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4404 a_411216_644902# mpw5_submission_0/isource_0/VM22D mpw5_submission_0/eigth_mirror_0/I_In vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4405 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4406 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4407 a_440818_643680# mpw5_submission_0/cmirror_channel_0/I_in_channel vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4408 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4409 mpw5_submission_0/outd_0/InputSignal io_analog[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4410 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4411 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4412 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4413 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4414 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4415 io_analog[1] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4416 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4417 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4418 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4419 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4420 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_434420_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4421 a_189936_651879# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4422 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4423 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4424 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4425 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4426 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4427 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4428 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4429 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4430 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4431 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4432 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4433 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4434 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4435 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4436 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4437 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4438 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_431720_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4439 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4440 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4441 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4442 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4443 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4444 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4445 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4446 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4447 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_184770_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4448 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4449 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4450 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4451 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4452 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4453 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4454 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4455 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4456 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4457 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4458 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4459 io_analog[6] mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/tia_core_0/Out_2 io_analog[6] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4460 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4461 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4462 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4463 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4464 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4465 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4466 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4467 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4468 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4469 vccd1 mpw5_submission_0/isource_0/VM14D mpw5_submission_0/isource_0/VM12G mpw5_submission_0/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4470 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4471 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4472 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4473 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4474 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4475 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4476 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4477 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4478 vssd1 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4479 vssd1 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4480 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_188820_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4481 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4482 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4483 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4484 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4485 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4486 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4487 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4488 mpw5_submission_0/tia_core_0/VM36D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM39D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4489 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4490 a_189936_651879# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4491 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4492 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4493 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_427670_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4494 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4495 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4496 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4497 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4498 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4499 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4500 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4501 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4502 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_186120_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4503 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4504 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4505 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4506 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4507 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4508 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4509 a_203370_649243# a_201520_649146# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4510 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4511 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4512 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4513 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4514 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4515 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4516 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4517 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4518 a_441658_643680# mpw5_submission_0/cmirror_channel_0/I_in_channel a_441720_645346# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4519 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4520 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4521 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4522 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4523 a_422158_661070# mpw5_submission_0/isource_0/VM11D vssd1 vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X4524 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4525 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4526 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4527 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4528 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4529 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4530 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4531 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4532 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4533 mpw5_submission_0/outd_0/V_da1_N vccd1 vssd1 sky130_fd_pr__res_high_po_2p85 l=6e+06u
X4534 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4535 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4536 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4537 a_190170_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4538 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4539 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4540 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4541 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4542 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/InputRef mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4543 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4544 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4545 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4546 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4547 mpw5_submission_0/outd_0/InputSignal io_analog[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4548 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4549 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4550 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4551 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4552 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4553 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4554 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4555 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4556 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4557 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4558 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4559 mpw5_submission_1/isource_0/VM3D mpw5_submission_1/isource_0/VM3G vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4560 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4561 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4562 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4563 mpw5_submission_0/outd_0/InputSignal io_analog[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4564 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4565 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4566 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4567 mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4568 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4569 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4570 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4571 vccd1 vssd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4572 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4573 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4574 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4575 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4576 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4577 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4578 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4579 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4580 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4581 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4582 mpw5_submission_1/outd_0/InputSignal io_analog[6] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4583 a_411216_644902# mpw5_submission_0/isource_0/VM22D mpw5_submission_0/eigth_mirror_0/I_In vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4584 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4585 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4586 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4587 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4588 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4589 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4590 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4591 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4592 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4593 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4594 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4595 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4596 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4597 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4598 mpw5_submission_1/isource_0/VM12G mpw5_submission_1/isource_0/VM14D vccd1 mpw5_submission_1/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4599 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4600 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4601 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4602 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4603 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4604 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4605 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4606 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4607 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4608 io_analog[0] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4609 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4610 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4611 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4612 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4613 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4614 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4615 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4616 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4617 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4618 a_200618_647480# mpw5_submission_1/cmirror_channel_0/I_in_channel vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4619 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4620 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4621 mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4622 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4623 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4624 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4625 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4626 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4627 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4628 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4629 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4630 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4631 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4632 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4633 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4634 mpw5_submission_0/eigth_mirror_0/I_out_5 mpw5_submission_0/eigth_mirror_0/I_In a_427670_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4635 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4636 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4637 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4638 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4639 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4640 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4641 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4642 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4643 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4644 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4645 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4646 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4647 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4648 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4649 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4650 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4651 a_431720_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4652 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4653 io_analog[6] mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/tia_core_0/Out_2 io_analog[6] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4654 vssd1 vccd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4655 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4656 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4657 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4658 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4659 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4660 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4661 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4662 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4663 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4664 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4665 vccd1 io_analog[1] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4666 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4667 a_434420_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4668 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4669 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4670 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4671 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4672 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4673 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4674 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4675 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4676 io_analog[0] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4677 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4678 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4679 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4680 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4681 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4682 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4683 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4684 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4685 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4686 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4687 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4688 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4689 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4690 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4691 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4692 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4693 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4694 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4695 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4696 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4697 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4698 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4699 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4700 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4701 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4702 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4703 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4704 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4705 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4706 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4707 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4708 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4709 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4710 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4711 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4712 mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4713 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4714 a_443850_641883# a_441720_645346# mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4715 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4716 mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/InputRef mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4717 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4718 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4719 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4720 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4721 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4722 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4723 a_433070_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4724 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4725 mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4726 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4727 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4728 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4729 a_186120_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4730 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4731 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4732 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4733 vssd1 vccd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4734 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4735 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4736 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4737 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4738 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4739 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4740 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4741 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4742 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4743 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4744 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4745 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4746 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4747 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4748 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4749 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4750 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4751 vssd1 io_analog[7] mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4752 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4753 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4754 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM36D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4755 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4756 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4757 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4758 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4759 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4760 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4761 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4762 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4763 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4764 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4765 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4766 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4767 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4768 mpw5_submission_0/tia_core_0/Out_2 mpw5_submission_0/outd_0/InputSignal io_analog[3] io_analog[3] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4769 vccd1 io_analog[1] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4770 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4771 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4772 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4773 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4774 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4775 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4776 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4777 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4778 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4779 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4780 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4781 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4782 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4783 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4784 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4785 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4786 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4787 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4788 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4789 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4790 a_203370_649243# a_201520_649146# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4791 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4792 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4793 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4794 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4795 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4796 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4797 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4798 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4799 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4800 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4801 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4802 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4803 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4804 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4805 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4806 a_443570_645443# a_441720_645346# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4807 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4808 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4809 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4810 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4811 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4812 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4813 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4814 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4815 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4816 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4817 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4818 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4819 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4820 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4821 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4822 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4823 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D36 vssd1 io_analog[3] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X4824 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4825 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4826 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_464438_656600# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4827 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4828 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4829 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4830 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4831 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4832 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4833 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4834 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4835 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4836 vssd1 mpw5_submission_0/isource_0/VM11D a_422158_661070# vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X4837 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4838 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4839 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4840 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4841 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4842 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4843 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4844 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4845 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4846 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4847 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4848 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4849 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4850 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4851 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4852 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4853 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4854 vccd1 io_analog[1] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4855 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4856 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4857 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4858 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4859 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4860 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4861 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4862 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4863 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4864 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4865 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4866 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4867 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4868 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4869 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4870 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4871 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4872 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4873 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4874 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4875 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4876 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4877 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4878 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4879 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4880 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4881 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4882 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4883 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4884 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4885 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4886 mpw5_submission_1/eigth_mirror_0/I_out_3 mpw5_submission_1/eigth_mirror_0/I_In a_190170_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4887 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4888 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4889 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4890 a_203650_645683# a_201520_649146# mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4891 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4892 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4893 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4894 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4895 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4896 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4897 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4898 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4899 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4900 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4901 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4902 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4903 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4904 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D37 io_analog[8] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X4905 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4906 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4907 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4908 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4909 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4910 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4911 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4912 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4913 a_434420_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4914 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4915 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4916 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4917 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4918 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4919 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4920 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4921 vccd1 io_analog[4] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4922 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4923 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4924 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4925 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4926 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4927 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4928 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4929 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4930 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4931 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4932 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4933 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4934 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4935 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4936 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4937 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4938 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4939 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4940 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4941 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4942 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4943 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4944 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4945 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4946 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4947 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4948 mpw5_submission_0/tia_core_0/VM5D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 io_analog[3] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4949 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4950 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4951 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4952 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4953 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4954 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4955 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4956 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4957 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4958 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4959 a_191520_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4960 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4961 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4962 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4963 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4964 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4965 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4966 a_201720_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4967 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4968 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4969 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4970 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4971 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4972 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4973 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4974 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4975 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4976 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4977 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4978 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4979 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4980 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4981 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4982 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4983 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4984 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4985 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4986 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4987 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4988 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4989 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4990 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4991 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4992 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4993 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4994 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4995 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4996 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4997 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4998 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4999 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5000 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5001 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5002 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5003 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5004 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5005 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5006 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5007 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5008 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5009 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5010 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5011 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5012 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5013 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5014 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5015 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5016 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5017 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5018 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5019 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5020 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5021 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5022 a_202298_647480# mpw5_submission_1/cmirror_channel_0/I_in_channel vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5023 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5024 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5025 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5026 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5027 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5028 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5029 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5030 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5031 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5032 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5033 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5034 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5035 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5036 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5037 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5038 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5039 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5040 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5041 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5042 io_analog[6] mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM5D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5043 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5044 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5045 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5046 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5047 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5048 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5049 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5050 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5051 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5052 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5053 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5054 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5055 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5056 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5057 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5058 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5059 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5060 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5061 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5062 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5063 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5064 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5065 mpw5_submission_0/eigth_mirror_0/I_out_2 mpw5_submission_0/eigth_mirror_0/I_In a_431720_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5066 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5067 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5068 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5069 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5070 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5071 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5072 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5073 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5074 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5075 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5076 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5077 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5078 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5079 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5080 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5081 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5082 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5083 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5084 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5085 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5086 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5087 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5088 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5089 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5090 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5091 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5092 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5093 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5094 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5095 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5096 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5097 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5098 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5099 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5100 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5101 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5102 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5103 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5104 mpw5_submission_1/tia_core_0/VM5D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5105 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5106 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5107 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5108 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5109 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5110 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5111 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5112 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5113 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5114 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5115 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5116 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5117 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5118 io_analog[3] mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/tia_core_0/Out_2 io_analog[3] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5119 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5120 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5121 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5122 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5123 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5124 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5125 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5126 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_424970_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5127 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5128 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5129 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5130 mpw5_submission_1/isource_0/VM3D a_171016_648702# mpw5_submission_1/isource_0/VM22D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X5131 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5132 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5133 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5134 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5135 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5136 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5137 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5138 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5139 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_427670_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5140 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5141 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5142 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5143 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5144 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5145 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5146 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5147 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5148 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5149 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5150 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5151 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5152 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5153 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5154 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5155 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5156 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5157 a_192870_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5158 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5159 mpw5_submission_0/tia_core_0/VM5D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 io_analog[3] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5160 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5161 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5162 io_analog[6] mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM5D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5163 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5164 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5165 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5166 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5167 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5168 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5169 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5170 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5171 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5172 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5173 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5174 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5175 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5176 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5177 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5178 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5179 mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5180 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5181 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5182 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5183 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5184 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5185 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5186 mpw5_submission_0/eigth_mirror_0/I_In mpw5_submission_0/isource_0/VM22D a_411216_644902# vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5187 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5188 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5189 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_426320_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5190 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5191 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5192 a_430136_648079# mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM14D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X5193 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5194 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5195 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5196 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5197 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5198 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5199 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5200 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_429020_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5201 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5202 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5203 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_426320_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5204 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5205 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5206 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5207 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5208 vssd1 mpw5_submission_1/cmirror_channel_0/I_in_channel a_201458_647480# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5209 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5210 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5211 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5212 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5213 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5214 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5215 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5216 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5217 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5218 a_203650_645683# a_201520_649146# mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
D38 vssd1 io_analog[3] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X5219 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5220 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5221 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5222 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5223 mpw5_submission_1/isource_0/VM8D a_181958_664870# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X5224 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5225 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5226 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5227 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5228 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5229 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5230 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5231 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5232 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5233 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5234 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5235 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5236 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5237 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5238 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5239 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5240 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5241 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5242 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5243 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5244 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5245 a_194220_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5246 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5247 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5248 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5249 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5250 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5251 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5252 vssd1 vccd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5253 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5254 mpw5_submission_1/outd_0/InputSignal io_analog[6] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5255 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5256 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5257 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5258 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5259 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5260 mpw5_submission_0/isource_0/VM12G mpw5_submission_0/isource_0/VM14D vccd1 mpw5_submission_0/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5261 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5262 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5263 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5264 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5265 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5266 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5267 a_430136_648079# mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM14D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X5268 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5269 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5270 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5271 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5272 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5273 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5274 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5275 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5276 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM36D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5277 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5278 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5279 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5280 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5281 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5282 a_181958_664870# mpw5_submission_1/isource_0/VM11D vssd1 vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X5283 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5284 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5285 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5286 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5287 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5288 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5289 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5290 a_189936_658659# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5291 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5292 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5293 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5294 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5295 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5296 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5297 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5298 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5299 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5300 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5301 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5302 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5303 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5304 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5305 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5306 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5307 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5308 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5309 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5310 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5311 vssd1 mpw5_submission_0/isource_0/VM12G mpw5_submission_0/isource_0/VM14D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X5312 vssd1 a_191036_648728# vssd1 sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X5313 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5314 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5315 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D39 vssd1 io_analog[3] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X5316 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5317 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5318 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5319 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5320 mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/InputRef mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5321 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5322 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5323 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5324 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5325 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5326 mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5327 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5328 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5329 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5330 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5331 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5332 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5333 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5334 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5335 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5336 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5337 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5338 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5339 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5340 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5341 a_191520_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5342 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5343 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5344 io_analog[6] mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM5D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5345 vccd1 io_analog[0] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5346 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5347 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5348 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5349 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5350 vssd1 mpw5_submission_1/cmirror_channel_0/I_in_channel a_202298_647480# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5351 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5352 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5353 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5354 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5355 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5356 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5357 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5358 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5359 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5360 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5361 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5362 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5363 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5364 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5365 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5366 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5367 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5368 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5369 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5370 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5371 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5372 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_654859# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5373 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5374 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5375 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5376 io_analog[0] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5377 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5378 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5379 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5380 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5381 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5382 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5383 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X5384 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5385 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5386 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5387 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5388 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5389 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5390 a_430136_654859# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5391 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5392 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5393 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5394 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5395 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5396 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5397 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5398 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5399 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5400 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5401 mpw5_submission_0/tia_core_0/VM36D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5402 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5403 mpw5_submission_1/isource_0/VM22D a_171016_648702# mpw5_submission_1/isource_0/VM3D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X5404 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5405 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5406 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5407 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5408 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5409 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5410 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5411 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5412 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5413 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5414 vccd1 a_441720_645346# a_441920_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5415 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5416 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5417 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5418 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5419 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5420 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5421 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5422 a_186120_640623# mpw5_submission_1/eigth_mirror_0/I_In mpw5_submission_1/eigth_mirror_0/I_out_6 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5423 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5424 vccd1 mpw5_submission_1/outd_0/V_da2_N vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5425 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5426 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5427 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5428 vssd1 mpw5_submission_0/cmirror_channel_0/I_in_channel a_440818_643680# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5429 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_431720_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5430 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5431 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5432 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5433 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5434 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5435 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5436 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5437 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5438 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5439 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5440 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_184770_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5441 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5442 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5443 a_429020_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5444 a_189936_651879# mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM14D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X5445 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5446 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5447 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5448 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5449 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5450 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5451 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5452 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5453 mpw5_submission_0/tia_core_0/VM6D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5454 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5455 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5456 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5457 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5458 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5459 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5460 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5461 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5462 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5463 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5464 mpw5_submission_1/eigth_mirror_0/I_out_2 mpw5_submission_1/eigth_mirror_0/I_In a_191520_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5465 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5466 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5467 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5468 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5469 mpw5_submission_1/outd_0/InputSignal io_analog[6] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5470 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5471 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5472 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5473 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5474 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5475 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5476 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5477 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5478 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5479 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5480 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5481 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5482 a_201720_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5483 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5484 mpw5_submission_0/eigth_mirror_0/I_In mpw5_submission_0/isource_0/VM22D a_411216_644902# vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5485 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5486 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5487 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5488 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5489 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5490 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5491 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5492 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5493 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5494 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_186120_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5495 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5496 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5497 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5498 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5499 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5500 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5501 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5502 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5503 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5504 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5505 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5506 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5507 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5508 a_189936_651879# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5509 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5510 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5511 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5512 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5513 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5514 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5515 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5516 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5517 mpw5_submission_0/outd_0/InputSignal io_analog[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5518 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D40 vssd1 io_analog[2] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X5519 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/InputRef mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5520 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5521 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5522 a_203370_649243# a_201520_649146# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5523 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5524 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5525 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5526 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5527 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5528 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5529 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5530 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5531 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5532 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5533 mpw5_submission_0/isource_0/VM14D mpw5_submission_0/isource_0/VM12G vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X5534 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5535 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5536 a_201520_649146# mpw5_submission_1/cmirror_channel_0/I_in_channel a_201458_647480# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5537 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5538 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5539 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5540 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5541 mpw5_submission_0/outd_0/InputSignal io_analog[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5542 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_649609# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5543 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5544 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5545 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5546 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5547 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5548 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5549 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5550 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5551 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5552 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5553 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5554 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5555 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5556 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5557 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5558 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5559 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5560 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5561 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5562 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5563 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5564 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5565 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5566 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
D41 vssd1 io_analog[0] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X5567 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X5568 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5569 a_433070_636823# mpw5_submission_0/eigth_mirror_0/I_In io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.74e+12p ps=1.374e+07u w=2e+06u l=200000u
X5570 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5571 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5572 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5573 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5574 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5575 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5576 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5577 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5578 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5579 a_189936_651879# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5580 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5581 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5582 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5583 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5584 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5585 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5586 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5587 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5588 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5589 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5590 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5591 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5592 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5593 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5594 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5595 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5596 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM31D mpw5_submission_0/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5597 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5598 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5599 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D42 vssd1 io_analog[8] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X5600 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5601 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5602 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5603 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5604 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5605 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5606 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5607 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5608 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5609 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5610 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5611 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5612 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5613 vssd1 mpw5_submission_1/isource_0/VM11D a_181958_664870# vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X5614 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5615 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5616 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5617 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5618 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5619 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5620 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5621 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5622 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5623 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5624 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5625 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5626 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5627 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5628 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5629 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5630 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5631 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5632 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5633 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5634 mpw5_submission_1/isource_0/VM3D a_171016_648702# mpw5_submission_1/isource_0/VM22D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X5635 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5636 mpw5_submission_1/isource_0/VM3D a_171016_648702# mpw5_submission_1/isource_0/VM22D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X5637 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5638 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5639 mpw5_submission_1/tia_core_0/Out_2 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5640 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5641 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5642 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5643 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5644 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5645 mpw5_submission_1/outd_0/InputSignal io_analog[6] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5646 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5647 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5648 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5649 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5650 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5651 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5652 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5653 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5654 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5655 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5656 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5657 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5658 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5659 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5660 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5661 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5662 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5663 vccd1 io_analog[1] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5664 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5665 a_422158_661070# mpw5_submission_0/isource_0/VM11D vssd1 vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X5666 a_184770_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5667 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5668 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5669 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5670 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5671 a_195570_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5672 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5673 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5674 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5675 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5676 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5677 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5678 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5679 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5680 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5681 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5682 a_434420_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5683 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5684 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X5685 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5686 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5687 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5688 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5689 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5690 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X5691 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5692 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5693 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5694 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5695 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5696 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5697 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5698 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5699 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5700 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5701 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5702 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5703 io_analog[3] mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/tia_core_0/Out_2 io_analog[3] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5704 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5705 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5706 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5707 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5708 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5709 vssd1 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X5710 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5711 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5712 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5713 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5714 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5715 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X5716 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5717 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5718 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5719 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5720 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5721 mpw5_submission_1/isource_0/VM12G a_184186_655038# vssd1 sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X5722 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5723 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5724 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
D43 vssd1 io_analog[1] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X5725 mpw5_submission_1/outd_0/InputSignal io_analog[6] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5726 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5727 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5728 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5729 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5730 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5731 mpw5_submission_0/tia_core_0/Out_2 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5732 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D44 io_analog[7] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X5733 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5734 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5735 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5736 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5737 a_433070_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5738 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5739 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5740 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5741 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5742 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5743 a_186120_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5744 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5745 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5746 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5747 io_analog[5] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5748 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5749 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5750 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5751 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5752 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5753 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5754 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5755 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5756 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5757 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5758 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5759 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5760 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5761 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5762 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5763 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5764 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5765 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5766 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5767 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5768 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5769 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5770 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5771 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5772 mpw5_submission_0/eigth_mirror_0/I_out_5 mpw5_submission_0/eigth_mirror_0/I_In a_427670_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5773 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5774 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5775 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5776 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5777 mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/InputRef mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5778 a_431720_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5779 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5780 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5781 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5782 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5783 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5784 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5785 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5786 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5787 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5788 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5789 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5790 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5791 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5792 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5793 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
D45 io_analog[3] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X5794 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5795 vssd1 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X5796 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5797 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5798 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5799 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5800 io_analog[6] mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/tia_core_0/Out_2 io_analog[6] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5801 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5802 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5803 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5804 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5805 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5806 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5807 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5808 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5809 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5810 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5811 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5812 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5813 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5814 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5815 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5816 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5817 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5818 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5819 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5820 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5821 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5822 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5823 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X5824 mpw5_submission_0/eigth_mirror_0/I_out_6 mpw5_submission_0/eigth_mirror_0/I_In a_426320_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5825 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5826 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5827 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5828 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5829 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5830 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5831 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5832 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5833 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5834 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5835 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5836 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5837 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5838 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5839 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5840 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5841 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5842 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5843 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5844 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5845 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5846 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5847 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5848 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5849 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5850 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5851 a_443850_641883# a_441720_645346# mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5852 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5853 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5854 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5855 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5856 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5857 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5858 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5859 a_188820_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5860 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5861 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5862 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5863 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5864 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5865 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5866 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5867 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5868 a_440818_643680# mpw5_submission_0/cmirror_channel_0/I_in_channel vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5869 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5870 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5871 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5872 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5873 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5874 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5875 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5876 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5877 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5878 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5879 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5880 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5881 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5882 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5883 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5884 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5885 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5886 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5887 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5888 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5889 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5890 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5891 mpw5_submission_1/tia_core_0/Out_2 mpw5_submission_1/outd_0/InputSignal io_analog[6] io_analog[6] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5892 vccd1 mpw5_submission_0/outd_0/V_da2_P vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5893 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5894 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5895 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5896 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5897 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5898 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5899 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5900 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5901 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5902 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5903 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5904 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5905 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5906 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5907 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5908 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5909 io_analog[5] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5910 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5911 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5912 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5913 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5914 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5915 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5916 vssd1 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X5917 vssd1 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X5918 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5919 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5920 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5921 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5922 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5923 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5924 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5925 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5926 io_analog[3] mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/tia_core_0/Out_2 io_analog[3] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5927 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5928 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5929 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5930 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5931 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5932 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5933 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5934 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5935 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5936 a_187470_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5937 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5938 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5939 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5940 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5941 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X5942 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5943 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5944 vccd1 io_analog[1] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5945 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5946 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
R1 vssd1 io_clamp_low[2] sky130_fd_pr__res_generic_m3 w=1.1e+07u l=250000u
X5947 mpw5_submission_0/tia_core_0/Out_2 mpw5_submission_0/outd_0/InputSignal io_analog[3] io_analog[3] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5948 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5949 a_441920_645443# a_441720_645346# a_441720_645346# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5950 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5951 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5952 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_192870_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5953 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5954 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5955 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5956 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5957 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5958 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5959 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5960 io_analog[5] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5961 io_analog[3] mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM5D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5962 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5963 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5964 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5965 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5966 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5967 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5968 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5969 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5970 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5971 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X5972 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5973 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5974 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5975 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5976 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5977 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5978 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5979 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5980 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5981 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5982 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5983 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5984 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5985 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5986 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5987 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5988 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5989 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5990 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5991 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5992 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5993 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5994 mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/InputRef mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5995 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5996 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D46 vssd1 io_analog[0] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X5997 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5998 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5999 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6000 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6001 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6002 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6003 vssd1 mpw5_submission_0/isource_0/VM11D a_422158_661070# vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X6004 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6005 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6006 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6007 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6008 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6009 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6010 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6011 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6012 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6013 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6014 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6015 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6016 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6017 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6018 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6019 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6020 vccd1 mpw5_submission_1/isource_0/VM14D mpw5_submission_1/isource_0/VM12G mpw5_submission_1/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6021 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6022 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6023 io_analog[3] mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/tia_core_0/Out_2 io_analog[3] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6024 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6025 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6026 vssd1 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6027 vssd1 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6028 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6029 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6030 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6031 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6032 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6033 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6034 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6035 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6036 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6037 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6038 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6039 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6040 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6041 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6042 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6043 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6044 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6045 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6046 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6047 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6048 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6049 vccd1 io_analog[0] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X6050 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6051 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6052 a_434420_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6053 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6054 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6055 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6056 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6057 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6058 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6059 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6060 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6061 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6062 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6063 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6064 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6065 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6066 vssd1 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM6D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6067 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6068 mpw5_submission_0/tia_core_0/VM36D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM39D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6069 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6070 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM31D mpw5_submission_1/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6071 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6072 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6073 a_430136_657119# mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM9D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X6074 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6075 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6076 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6077 a_431720_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6078 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6079 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6080 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6081 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6082 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6083 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6084 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6085 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6086 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D47 io_analog[8] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X6087 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6088 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6089 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6090 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6091 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6092 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6093 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6094 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6095 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6096 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6097 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6098 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6099 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6100 mpw5_submission_1/outd_0/V_da1_N vccd1 vssd1 sky130_fd_pr__res_high_po_2p85 l=6e+06u
X6101 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6102 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6103 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6104 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6105 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6106 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6107 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6108 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6109 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6110 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6111 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6112 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6113 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6114 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6115 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6116 io_analog[6] mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/tia_core_0/Out_2 io_analog[6] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6117 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6118 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6119 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6120 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6121 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6122 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6123 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_188820_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6124 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6125 a_430370_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6126 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6127 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6128 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6129 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6130 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6131 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6132 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6133 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6134 mpw5_submission_1/tia_core_0/VM5D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 io_analog[6] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6135 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6136 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6137 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6138 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6139 a_189936_651879# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6140 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6141 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6142 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_427670_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6143 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6144 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6145 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6146 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6147 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6148 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6149 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6150 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6151 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6152 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6153 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6154 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6155 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6156 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6157 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6158 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6159 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6160 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6161 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6162 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6163 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6164 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6165 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6166 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6167 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6168 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6169 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6170 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6171 vssd1 vccd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
D48 vssd1 io_analog[0] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X6172 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6173 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6174 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6175 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6176 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6177 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6178 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6179 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6180 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6181 mpw5_submission_1/eigth_mirror_0/I_out_5 mpw5_submission_1/eigth_mirror_0/I_In a_187470_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6182 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6183 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6184 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6185 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6186 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6187 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6188 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6189 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6190 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6191 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6192 io_analog[4] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X6193 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6194 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6195 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6196 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6197 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224238_660400# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6198 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6199 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6200 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6201 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6202 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6203 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_429020_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6204 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6205 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6206 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6207 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_426320_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6208 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6209 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6210 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6211 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6212 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6213 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6214 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6215 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6216 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6217 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6218 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6219 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6220 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6221 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6222 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6223 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6224 vccd1 io_analog[5] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X6225 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6226 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6227 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6228 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6229 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6230 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6231 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6232 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6233 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6234 mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__cap_var_lvt pd=0u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X6235 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6236 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6237 io_analog[4] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X6238 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6239 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6240 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6241 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6242 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6243 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6244 mpw5_submission_1/eigth_mirror_0/I_out_6 mpw5_submission_1/eigth_mirror_0/I_In a_186120_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6245 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6246 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6247 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6248 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6249 mpw5_submission_0/tia_core_0/Out_2 mpw5_submission_0/outd_0/InputSignal io_analog[3] io_analog[3] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6250 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6251 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6252 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_424970_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6253 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6254 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6255 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6256 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6257 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6258 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6259 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6260 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6261 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6262 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6263 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6264 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6265 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6266 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6267 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6268 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6269 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6270 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6271 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6272 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6273 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6274 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6275 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6276 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6277 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6278 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6279 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6280 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6281 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6282 a_430136_648079# mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM14D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X6283 a_411216_644902# mpw5_submission_0/isource_0/VM22D mpw5_submission_0/eigth_mirror_0/I_In vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6284 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM31D mpw5_submission_1/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6285 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6286 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6287 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6288 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6289 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6290 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6291 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6292 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6293 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6294 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6295 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6296 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6297 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6298 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6299 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6300 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6301 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6302 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6303 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6304 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6305 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6306 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6307 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6308 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6309 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6310 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6311 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6312 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6313 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6314 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6315 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_426320_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6316 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6317 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6318 mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/InputRef mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6319 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6320 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6321 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6322 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6323 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6324 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6325 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6326 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6327 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6328 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6329 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6330 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6331 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6332 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6333 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6334 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6335 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6336 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6337 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6338 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6339 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6340 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6341 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6342 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6343 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6344 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6345 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6346 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6347 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6348 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6349 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6350 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6351 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6352 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6353 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6354 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6355 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6356 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6357 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6358 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6359 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6360 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6361 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6362 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6363 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6364 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6365 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6366 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6367 a_430136_648079# mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM14D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X6368 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6369 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6370 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6371 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6372 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6373 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6374 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6375 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6376 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6377 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6378 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6379 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6380 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6381 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6382 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6383 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6384 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6385 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6386 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6387 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6388 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6389 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6390 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6391 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6392 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6393 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6394 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6395 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6396 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6397 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6398 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6399 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6400 mpw5_submission_0/tia_core_0/VM6D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6401 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6402 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6403 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6404 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6405 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6406 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6407 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6408 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6409 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6410 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6411 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6412 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6413 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6414 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6415 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6416 a_203370_649243# a_201520_649146# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6417 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6418 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6419 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6420 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6421 mpw5_submission_0/tia_core_0/VM31D mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6422 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6423 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6424 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6425 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6426 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6427 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6428 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/InputRef mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6429 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6430 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6431 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6432 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6433 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6434 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6435 a_181958_664870# mpw5_submission_1/isource_0/VM11D vssd1 vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X6436 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6437 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6438 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6439 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6440 a_190170_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6441 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6442 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6443 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6444 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6445 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6446 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6447 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6448 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D49 vssd1 io_analog[3] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X6449 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6450 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6451 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6452 a_429020_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6453 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6454 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6455 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6456 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6457 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6458 a_187470_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6459 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6460 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6461 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6462 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6463 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6464 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6465 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6466 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6467 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6468 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6469 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6470 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6471 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6472 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6473 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6474 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6475 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6476 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6477 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6478 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6479 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6480 vccd1 mpw5_submission_1/outd_0/V_da2_N vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X6481 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6482 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6483 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6484 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6485 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6486 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6487 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6488 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6489 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6490 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6491 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6492 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6493 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6494 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6495 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6496 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6497 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6498 vccd1 io_analog[4] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X6499 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6500 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6501 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6502 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6503 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6504 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6505 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6506 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6507 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6508 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6509 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6510 mpw5_submission_0/eigth_mirror_0/I_In mpw5_submission_0/isource_0/VM22D a_411216_644902# vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6511 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6512 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6513 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6514 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6515 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6516 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6517 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6518 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6519 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6520 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6521 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6522 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6523 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6524 a_422158_661070# mpw5_submission_0/isource_0/VM11D vssd1 vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X6525 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6526 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6527 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6528 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6529 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6530 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6531 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6532 vccd1 vssd1 mpw5_submission_1/tia_core_0/VM31D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6533 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6534 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6535 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6536 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6537 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6538 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6539 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6540 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6541 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6542 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6543 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6544 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6545 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6546 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6547 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6548 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6549 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6550 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6551 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6552 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6553 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6554 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6555 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6556 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6557 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6558 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6559 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6560 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6561 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6562 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D50 io_analog[1] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X6563 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/InputRef mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6564 mpw5_submission_0/outd_0/InputSignal io_analog[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6565 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6566 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6567 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6568 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6569 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D51 vssd1 io_analog[0] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X6570 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6571 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6572 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6573 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6574 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6575 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6576 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6577 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6578 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6579 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6580 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6581 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6582 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6583 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6584 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6585 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6586 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6587 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6588 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6589 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6590 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6591 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6592 mpw5_submission_1/eigth_mirror_0/I_out_2 mpw5_submission_1/eigth_mirror_0/I_In a_191520_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6593 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6594 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6595 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6596 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6597 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6598 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6599 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6600 mpw5_submission_1/outd_0/InputSignal io_analog[6] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6601 mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__cap_var_lvt pd=0u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X6602 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6603 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6604 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
R2 vssd1 io_clamp_low[0] sky130_fd_pr__res_generic_m3 w=1.1e+07u l=250000u
X6605 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6606 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6607 a_443850_641883# a_441720_645346# mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6608 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6609 mpw5_submission_1/eigth_mirror_0/I_In mpw5_submission_1/isource_0/VM22D a_171016_648702# vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6610 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6611 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6612 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6613 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6614 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6615 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6616 vccd1 vssd1 mpw5_submission_0/tia_core_0/VM31D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6617 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6618 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6619 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6620 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6621 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6622 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6623 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6624 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6625 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_435770_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6626 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6627 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6628 a_435770_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6629 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6630 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6631 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6632 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6633 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6634 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6635 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6636 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6637 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6638 a_203370_649243# a_201520_649146# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6639 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6640 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6641 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6642 vssd1 io_analog[7] mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6643 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6644 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6645 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6646 a_189936_651879# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6647 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6648 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6649 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6650 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6651 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6652 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6653 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6654 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6655 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6656 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6657 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6658 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6659 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6660 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6661 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6662 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6663 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6664 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6665 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6666 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6667 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6668 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6669 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6670 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6671 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6672 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6673 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6674 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6675 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6676 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6677 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6678 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6679 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6680 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6681 a_430136_645809# mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM22D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X6682 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6683 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6684 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6685 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6686 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6687 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6688 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6689 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6690 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6691 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6692 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6693 io_analog[6] mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/tia_core_0/Out_2 io_analog[6] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6694 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6695 a_430136_648079# mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM14D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X6696 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6697 a_441920_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6698 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6699 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6700 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6701 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6702 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6703 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6704 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6705 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6706 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6707 mpw5_submission_0/outd_0/V_da2_N vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X6708 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6709 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6710 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6711 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6712 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6713 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6714 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D52 io_analog[8] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X6715 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6716 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6717 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6718 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6719 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6720 mpw5_submission_1/tia_core_0/VM36D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6721 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6722 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6723 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6724 io_analog[0] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X6725 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6726 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6727 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6728 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6729 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6730 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM31D mpw5_submission_0/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6731 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6732 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6733 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6734 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6735 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6736 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6737 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6738 a_441720_645346# a_441720_645346# a_441920_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6739 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6740 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6741 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6742 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6743 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6744 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6745 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6746 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6747 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6748 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6749 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6750 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6751 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6752 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6753 vssd1 mpw5_submission_1/isource_0/VM11D a_181958_664870# vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X6754 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6755 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6756 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6757 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6758 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D53 io_analog[0] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X6759 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6760 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6761 vssd1 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6762 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6763 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6764 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6765 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6766 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6767 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6768 io_analog[5] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X6769 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6770 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/InputRef mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6771 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6772 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6773 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6774 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6775 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6776 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6777 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6778 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6779 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6780 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6781 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6782 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6783 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6784 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6785 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6786 mpw5_submission_1/outd_0/InputSignal io_analog[6] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6787 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6788 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6789 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6790 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6791 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6792 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6793 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6794 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6795 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6796 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6797 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_190170_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6798 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6799 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6800 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6801 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6802 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6803 mpw5_submission_1/isource_0/VM12G mpw5_submission_1/isource_0/VM14D vccd1 mpw5_submission_1/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6804 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6805 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6806 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6807 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6808 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6809 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6810 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6811 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6812 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6813 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6814 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6815 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D54 vssd1 io_analog[8] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X6816 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6817 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6818 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6819 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6820 mpw5_submission_0/tia_core_0/Out_2 mpw5_submission_0/outd_0/InputSignal io_analog[3] io_analog[3] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6821 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6822 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6823 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6824 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6825 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6826 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6827 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6828 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6829 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6830 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6831 a_426320_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6832 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6833 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6834 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6835 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6836 mpw5_submission_0/isource_0/VM3G a_425526_651238# vssd1 sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X6837 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6838 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6839 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6840 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6841 a_201458_647480# mpw5_submission_1/cmirror_channel_0/I_in_channel vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6842 a_443570_645443# a_441720_645346# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6843 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6844 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6845 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6846 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6847 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6848 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6849 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6850 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6851 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6852 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_191520_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6853 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6854 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6855 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6856 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6857 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6858 vssd1 mpw5_submission_1/isource_0/VM12G mpw5_submission_1/isource_0/VM14D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6859 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6860 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6861 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6862 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6863 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6864 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6865 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6866 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6867 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6868 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6869 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6870 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6871 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6872 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6873 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6874 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6875 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6876 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6877 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6878 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6879 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6880 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6881 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6882 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6883 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6884 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6885 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6886 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6887 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6888 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6889 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6890 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6891 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6892 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6893 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6894 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6895 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6896 vccd1 io_analog[4] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X6897 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6898 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6899 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_649609# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6900 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6901 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6902 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6903 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6904 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6905 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6906 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6907 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6908 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6909 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6910 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6911 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6912 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6913 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6914 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6915 mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__cap_var_lvt pd=0u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X6916 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6917 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6918 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6919 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6920 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6921 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6922 io_analog[4] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X6923 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_658659# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6924 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6925 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6926 io_analog[6] mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM5D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6927 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6928 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6929 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6930 a_429646_642496# a_411216_644902# vssd1 sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X6931 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6932 mpw5_submission_1/tia_core_0/Out_2 mpw5_submission_1/outd_0/InputSignal io_analog[6] io_analog[6] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6933 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6934 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6935 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6936 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6937 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6938 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6939 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_192870_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6940 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6941 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6942 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6943 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6944 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6945 a_189936_658659# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6946 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6947 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6948 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6949 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6950 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6951 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6952 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/Disable_TIA vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D55 io_analog[2] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X6953 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6954 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6955 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6956 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6957 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6958 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6959 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6960 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6961 mpw5_submission_1/isource_0/VM3D a_171016_648702# mpw5_submission_1/isource_0/VM22D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6962 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6963 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6964 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6965 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6966 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6967 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6968 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6969 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6970 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6971 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6972 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6973 a_435770_636823# mpw5_submission_0/eigth_mirror_0/I_In mpw5_submission_0/eigth_mirror_0/I_In vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6974 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6975 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6976 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6977 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6978 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6979 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6980 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6981 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6982 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6983 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6984 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6985 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6986 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6987 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6988 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6989 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6990 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6991 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6992 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6993 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6994 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6995 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6996 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6997 mpw5_submission_1/outd_0/V_da2_P vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X6998 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6999 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7000 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_657119# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7001 vssd1 mpw5_submission_1/cmirror_channel_0/I_in_channel a_200618_647480# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7002 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D56 io_analog[7] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X7003 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7004 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7005 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7006 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7007 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7008 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7009 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7010 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7011 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7012 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7013 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7014 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7015 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7016 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7017 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7018 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7019 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7020 a_434420_636823# mpw5_submission_0/eigth_mirror_0/I_In mpw5_submission_0/cmirror_channel_0/I_in_channel vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7021 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7022 mpw5_submission_1/tia_core_0/Out_2 mpw5_submission_1/outd_0/InputSignal io_analog[6] io_analog[6] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7023 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7024 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7025 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7026 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7027 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7028 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_654859# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7029 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7030 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7031 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7032 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7033 vssd1 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM36D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7034 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7035 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7036 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7037 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7038 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7039 io_analog[3] mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/tia_core_0/Out_2 io_analog[3] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7040 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7041 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7042 a_192870_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7043 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7044 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7045 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7046 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7047 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7048 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7049 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7050 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7051 a_431720_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7052 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7053 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7054 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7055 vccd1 a_441720_645346# a_441920_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7056 mpw5_submission_1/isource_0/VM14D mpw5_submission_1/isource_0/VM12G vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X7057 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7058 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7059 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7060 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7061 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7062 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7063 vccd1 io_analog[5] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X7064 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7065 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7066 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7067 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7068 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7069 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7070 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7071 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7072 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7073 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7074 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7075 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7076 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7077 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7078 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7079 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7080 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7081 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X7082 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7083 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7084 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7085 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7086 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7087 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7088 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7089 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7090 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7091 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7092 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7093 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7094 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7095 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7096 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7097 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7098 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7099 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7100 a_192870_640623# mpw5_submission_1/eigth_mirror_0/I_In mpw5_submission_1/eigth_mirror_0/I_out_1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7101 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7102 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7103 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7104 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7105 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7106 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7107 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7108 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7109 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7110 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7111 a_430370_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7112 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7113 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7114 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7115 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7116 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7117 mpw5_submission_0/isource_0/VM12G mpw5_submission_0/isource_0/VM14D vccd1 mpw5_submission_0/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7118 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7119 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7120 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7121 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7122 mpw5_submission_0/tia_core_0/Out_2 mpw5_submission_0/outd_0/InputSignal io_analog[3] io_analog[3] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7123 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7124 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7125 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7126 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7127 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7128 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7129 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7130 a_427670_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7131 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7132 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7133 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7134 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7135 a_443570_645443# a_441720_645346# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7136 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7137 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7138 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7139 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7140 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7141 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7142 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7143 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7144 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7145 io_analog[3] mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/tia_core_0/Out_2 io_analog[3] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7146 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7147 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7148 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7149 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7150 vssd1 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM36D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7151 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X7152 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7153 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7154 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7155 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7156 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7157 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7158 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7159 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7160 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7161 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7162 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7163 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7164 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7165 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7166 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7167 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7168 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7169 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7170 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7171 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7172 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7173 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7174 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7175 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7176 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7177 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7178 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7179 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7180 vccd1 a_441720_645346# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7181 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7182 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7183 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7184 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7185 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7186 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7187 mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/InputRef mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7188 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7189 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7190 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7191 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7192 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7193 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7194 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7195 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7196 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7197 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7198 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7199 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7200 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7201 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7202 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7203 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7204 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7205 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7206 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
D57 vssd1 io_analog[8] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X7207 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7208 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7209 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7210 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7211 a_189936_651879# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7212 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7213 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7214 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7215 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7216 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7217 vssd1 vccd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7218 vssd1 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X7219 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7220 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7221 vccd1 a_201520_649146# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7222 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7223 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7224 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7225 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7226 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7227 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D58 io_analog[8] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X7228 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7229 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7230 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7231 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7232 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7233 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7234 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7235 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7236 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7237 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7238 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X7239 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7240 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7241 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7242 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7243 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7244 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7245 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7246 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7247 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7248 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7249 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7250 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7251 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7252 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7253 a_434420_636823# mpw5_submission_0/eigth_mirror_0/I_In mpw5_submission_0/cmirror_channel_0/I_in_channel vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7254 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7255 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7256 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7257 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7258 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7259 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7260 a_202298_647480# mpw5_submission_1/cmirror_channel_0/I_in_channel vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7261 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7262 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7263 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D59 vssd1 io_analog[7] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X7264 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7265 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7266 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7267 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7268 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7269 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7270 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7271 io_analog[1] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X7272 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7273 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7274 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7275 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7276 mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__cap_var_lvt pd=0u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X7277 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7278 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7279 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7280 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7281 a_411216_644902# mpw5_submission_0/isource_0/VM22D mpw5_submission_0/eigth_mirror_0/I_In vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7282 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7283 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7284 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7285 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM31D mpw5_submission_0/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7286 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7287 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7288 a_443850_641883# a_441720_645346# mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7289 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7290 mpw5_submission_1/eigth_mirror_0/I_out_5 mpw5_submission_1/eigth_mirror_0/I_In a_187470_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7291 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7292 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7293 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7294 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7295 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7296 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7297 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7298 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7299 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7300 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7301 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7302 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7303 a_430136_648079# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7304 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7305 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7306 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7307 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7308 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7309 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7310 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7311 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7312 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7313 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7314 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7315 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7316 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7317 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7318 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7319 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7320 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7321 vssd1 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X7322 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7323 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7324 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7325 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7326 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7327 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7328 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7329 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7330 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7331 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7332 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7333 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7334 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7335 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7336 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7337 mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/InputRef mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7338 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7339 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7340 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7341 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7342 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7343 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7344 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7345 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7346 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7347 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7348 mpw5_submission_1/eigth_mirror_0/I_out_6 mpw5_submission_1/eigth_mirror_0/I_In a_186120_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7349 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7350 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X7351 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7352 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7353 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7354 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7355 vccd1 mpw5_submission_0/isource_0/VM14D mpw5_submission_0/isource_0/VM12G mpw5_submission_0/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7356 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7357 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7358 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7359 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7360 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7361 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7362 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7363 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7364 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7365 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/InputRef mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7366 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7367 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7368 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7369 a_442498_643680# mpw5_submission_0/cmirror_channel_0/I_in_channel vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7370 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7371 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7372 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7373 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7374 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7375 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7376 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7377 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7378 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7379 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7380 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7381 a_171016_648702# mpw5_submission_1/isource_0/VM22D mpw5_submission_1/eigth_mirror_0/I_In vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7382 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7383 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM31D mpw5_submission_1/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7384 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7385 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7386 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7387 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7388 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7389 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7390 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7391 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7392 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7393 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7394 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7395 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7396 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7397 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7398 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7399 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7400 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7401 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7402 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7403 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7404 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7405 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7406 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7407 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7408 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7409 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7410 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7411 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7412 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7413 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 io_analog[7] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7414 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7415 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7416 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7417 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7418 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7419 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7420 a_187470_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7421 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7422 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7423 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7424 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7425 vssd1 mpw5_submission_1/cmirror_channel_0/I_in_channel a_201458_647480# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7426 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7427 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7428 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7429 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7430 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7431 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7432 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7433 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7434 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7435 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7436 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7437 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7438 vccd1 io_analog[5] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X7439 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7440 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7441 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7442 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7443 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7444 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7445 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7446 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7447 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7448 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7449 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7450 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7451 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7452 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7453 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7454 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7455 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7456 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7457 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7458 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X7459 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7460 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7461 mpw5_submission_1/tia_core_0/VM31D mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7462 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7463 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7464 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7465 a_426056_648806# a_425526_651238# vssd1 sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X7466 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7467 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7468 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7469 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7470 mpw5_submission_1/tia_core_0/VM31D vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7471 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7472 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7473 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7474 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7475 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7476 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7477 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7478 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7479 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7480 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7481 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7482 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7483 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM31D mpw5_submission_0/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7484 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7485 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7486 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7487 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7488 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7489 io_analog[1] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X7490 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7491 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7492 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7493 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7494 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7495 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7496 a_189936_651879# mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM14D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X7497 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7498 a_189936_660919# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7499 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7500 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7501 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7502 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7503 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7504 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7505 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7506 mpw5_submission_0/tia_core_0/VM31D mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7507 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7508 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7509 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7510 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7511 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7512 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7513 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7514 mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/InputRef mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7515 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7516 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7517 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7518 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_187470_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7519 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7520 a_184770_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7521 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7522 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7523 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7524 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7525 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7526 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7527 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7528 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7529 vssd1 mpw5_submission_0/cmirror_channel_0/I_in_channel a_441658_643680# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7530 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7531 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7532 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7533 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7534 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7535 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7536 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7537 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7538 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7539 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7540 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7541 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_192870_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7542 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7543 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7544 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7545 vccd1 io_analog[4] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X7546 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7547 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7548 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7549 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X7550 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7551 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7552 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7553 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7554 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7555 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7556 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7557 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7558 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7559 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7560 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7561 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7562 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7563 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7564 a_171016_648702# mpw5_submission_1/isource_0/VM22D mpw5_submission_1/eigth_mirror_0/I_In vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7565 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7566 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7567 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7568 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7569 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7570 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7571 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7572 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7573 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7574 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7575 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X7576 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7577 a_189936_651879# mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM14D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X7578 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7579 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7580 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X7581 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7582 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7583 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7584 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM31D mpw5_submission_0/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7585 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7586 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7587 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7588 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7589 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7590 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7591 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7592 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_645809# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7593 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7594 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7595 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7596 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_435770_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7597 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7598 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7599 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7600 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7601 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7602 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7603 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7604 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X7605 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_194220_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7606 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7607 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7608 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7609 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7610 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7611 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7612 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7613 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7614 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7615 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7616 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7617 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7618 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7619 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7620 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7621 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7622 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7623 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7624 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7625 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7626 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7627 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7628 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7629 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7630 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7631 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7632 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7633 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7634 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7635 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7636 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7637 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7638 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7639 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7640 mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7641 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7642 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7643 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7644 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7645 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7646 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7647 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7648 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7649 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7650 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7651 vssd1 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM5D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7652 a_201720_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7653 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7654 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7655 vssd1 mpw5_submission_0/cmirror_channel_0/I_in_channel a_440818_643680# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7656 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7657 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7658 io_analog[0] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X7659 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7660 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7661 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7662 mpw5_submission_1/tia_core_0/VM6D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7663 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7664 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7665 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7666 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7667 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7668 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7669 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7670 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7671 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7672 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7673 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7674 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7675 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7676 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7677 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7678 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7679 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7680 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7681 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7682 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7683 io_analog[1] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X7684 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7685 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7686 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7687 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7688 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7689 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7690 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM31D mpw5_submission_1/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7691 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7692 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7693 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7694 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7695 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7696 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7697 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7698 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7699 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7700 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7701 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7702 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7703 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7704 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7705 a_189936_651879# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7706 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7707 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7708 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7709 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7710 mpw5_submission_1/outd_0/InputSignal io_analog[6] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7711 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7712 a_435770_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7713 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7714 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7715 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7716 a_201720_649243# a_201520_649146# a_201520_649146# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7717 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7718 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7719 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7720 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7721 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7722 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7723 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7724 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7725 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7726 a_188820_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7727 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_430370_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7728 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7729 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7730 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7731 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7732 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7733 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7734 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7735 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7736 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7737 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7738 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7739 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7740 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7741 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7742 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7743 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7744 mpw5_submission_0/eigth_mirror_0/I_In mpw5_submission_0/eigth_mirror_0/I_In a_435770_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7745 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7746 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7747 io_analog[0] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X7748 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7749 mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7750 a_430136_648079# mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM14D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X7751 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7752 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7753 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7754 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7755 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7756 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7757 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7758 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7759 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7760 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7761 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7762 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7763 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7764 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7765 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7766 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7767 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7768 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7769 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7770 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7771 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_658659# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7772 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7773 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7774 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7775 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7776 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7777 a_187470_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7778 mpw5_submission_1/tia_core_0/Out_2 mpw5_submission_1/outd_0/InputSignal io_analog[6] io_analog[6] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7779 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7780 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7781 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7782 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7783 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7784 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7785 vssd1 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X7786 vssd1 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X7787 a_426320_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7788 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7789 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7790 io_analog[6] mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/tia_core_0/Out_2 io_analog[6] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7791 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7792 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7793 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7794 a_184770_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7795 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7796 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7797 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7798 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7799 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7800 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7801 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7802 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7803 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7804 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D60 vssd1 io_analog[2] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X7805 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7806 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7807 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7808 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7809 mpw5_submission_0/tia_core_0/VM31D mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7810 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D61 io_analog[1] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X7811 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X7812 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7813 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7814 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7815 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7816 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7817 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7818 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7819 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7820 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7821 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7822 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7823 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7824 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7825 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7826 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7827 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7828 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7829 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7830 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7831 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7832 a_441720_645346# a_441720_645346# a_441920_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7833 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7834 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7835 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7836 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7837 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7838 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7839 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7840 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7841 a_464438_656600# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7842 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7843 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7844 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7845 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7846 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7847 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7848 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7849 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7850 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7851 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7852 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7853 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7854 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7855 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7856 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7857 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7858 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7859 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7860 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7861 mpw5_submission_1/isource_0/VM3D a_171016_648702# mpw5_submission_1/isource_0/VM22D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X7862 vccd1 vssd1 mpw5_submission_0/tia_core_0/VM31D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7863 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7864 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7865 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7866 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7867 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7868 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7869 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7870 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7871 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7872 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7873 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7874 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7875 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7876 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7877 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7878 vccd1 mpw5_submission_0/isource_0/VM14D mpw5_submission_0/isource_0/VM12G mpw5_submission_0/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7879 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7880 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7881 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7882 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7883 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7884 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7885 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7886 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7887 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7888 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7889 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7890 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7891 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7892 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7893 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7894 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7895 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7896 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7897 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7898 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7899 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7900 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7901 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7902 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7903 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7904 mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7905 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7906 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7907 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7908 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7909 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7910 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7911 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7912 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7913 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7914 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7915 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7916 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7917 a_443570_645443# a_441720_645346# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7918 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7919 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7920 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7921 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7922 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7923 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7924 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7925 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7926 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7927 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7928 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7929 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7930 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7931 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7932 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7933 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7934 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7935 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7936 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7937 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7938 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7939 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7940 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7941 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7942 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7943 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7944 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7945 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7946 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7947 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7948 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7949 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7950 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7951 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7952 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7953 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7954 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7955 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7956 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7957 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7958 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7959 io_analog[0] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X7960 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7961 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7962 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7963 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7964 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7965 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7966 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7967 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7968 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7969 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7970 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7971 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7972 vssd1 vccd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7973 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7974 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7975 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7976 a_443570_645443# a_441720_645346# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7977 a_443850_641883# a_441720_645346# mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7978 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7979 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7980 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7981 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7982 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7983 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7984 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7985 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7986 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7987 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7988 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7989 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7990 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7991 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7992 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7993 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7994 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7995 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7996 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7997 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7998 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7999 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8000 a_429020_636823# mpw5_submission_0/eigth_mirror_0/I_In mpw5_submission_0/eigth_mirror_0/I_out_4 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
D62 io_analog[0] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X8001 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8002 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8003 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8004 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8005 a_203650_645683# a_201520_649146# mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8006 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8007 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8008 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8009 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8010 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8011 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8012 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8013 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8014 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8015 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8016 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8017 mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8018 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8019 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8020 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8021 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8022 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8023 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8024 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8025 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8026 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8027 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8028 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8029 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8030 mpw5_submission_1/tia_core_0/Out_2 mpw5_submission_1/outd_0/InputSignal io_analog[6] io_analog[6] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8031 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8032 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8033 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8034 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8035 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8036 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8037 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8038 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8039 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8040 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8041 a_443850_641883# a_441720_645346# mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8042 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8043 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8044 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8045 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8046 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8047 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8048 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8049 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8050 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8051 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8052 a_440818_643680# mpw5_submission_0/cmirror_channel_0/I_in_channel mpw5_submission_0/cmirror_channel_0/I_in_channel vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8053 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8054 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8055 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8056 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8057 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8058 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8059 mpw5_submission_0/eigth_mirror_0/I_In mpw5_submission_0/isource_0/VM22D a_411216_644902# vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8060 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
D63 vssd1 io_analog[7] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X8061 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8062 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8063 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8064 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8065 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8066 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8067 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8068 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8069 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8070 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8071 a_203370_649243# a_201520_649146# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8072 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8073 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8074 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8075 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8076 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8077 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D64 io_analog[0] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X8078 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8079 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8080 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8081 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8082 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8083 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8084 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8085 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8086 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8087 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8088 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8089 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8090 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8091 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8092 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8093 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8094 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8095 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8096 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8097 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8098 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8099 mpw5_submission_1/isource_0/VM22D a_171016_648702# mpw5_submission_1/isource_0/VM3D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X8100 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8101 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8102 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8103 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8104 a_430136_657119# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8105 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8106 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8107 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8108 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8109 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8110 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8111 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8112 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8113 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8114 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8115 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8116 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/InputRef mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8117 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8118 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8119 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8120 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8121 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/InputRef mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8122 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8123 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8124 io_analog[6] mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/tia_core_0/Out_2 io_analog[6] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8125 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8126 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8127 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8128 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8129 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8130 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8131 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8132 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8133 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8134 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8135 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8136 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8137 mpw5_submission_0/isource_0/VM12G mpw5_submission_0/isource_0/VM14D vccd1 mpw5_submission_0/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8138 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8139 mpw5_submission_1/tia_core_0/Out_2 mpw5_submission_1/outd_0/InputSignal io_analog[6] io_analog[6] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8140 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8141 mpw5_submission_0/isource_0/VM12G mpw5_submission_0/isource_0/VM14D vccd1 mpw5_submission_0/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8142 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8143 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8144 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8145 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8146 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8147 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8148 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8149 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8150 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8151 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8152 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8153 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8154 mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/InputRef mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8155 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8156 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8157 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8158 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8159 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8160 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8161 vssd1 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X8162 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8163 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8164 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8165 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8166 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8167 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8168 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8169 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8170 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8171 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8172 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8173 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8174 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8175 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8176 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8177 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8178 mpw5_submission_1/eigth_mirror_0/I_In mpw5_submission_1/isource_0/VM22D a_171016_648702# vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8179 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8180 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8181 vccd1 vssd1 mpw5_submission_1/tia_core_0/VM31D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8182 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8183 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8184 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8185 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8186 io_analog[5] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X8187 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8188 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8189 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8190 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8191 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8192 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8193 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8194 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8195 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8196 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8197 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8198 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8199 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8200 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8201 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8202 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8203 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8204 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8205 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8206 vccd1 mpw5_submission_0/outd_0/V_da2_N vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X8207 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8208 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8209 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D65 io_analog[2] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X8210 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8211 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8212 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8213 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8214 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8215 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8216 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8217 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8218 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8219 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8220 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8221 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8222 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8223 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8224 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8225 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8226 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8227 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8228 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8229 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8230 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8231 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8232 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8233 a_427670_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8234 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8235 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8236 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8237 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8238 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8239 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8240 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8241 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8242 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8243 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_433070_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8244 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8245 mpw5_submission_0/tia_core_0/Out_2 mpw5_submission_0/outd_0/InputSignal io_analog[3] io_analog[3] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8246 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8247 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8248 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8249 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8250 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8251 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8252 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_435770_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8253 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8254 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8255 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8256 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8257 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8258 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8259 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8260 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8261 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8262 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8263 vssd1 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X8264 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8265 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8266 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X8267 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8268 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8269 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8270 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8271 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8272 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8273 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8274 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8275 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8276 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM31D mpw5_submission_1/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8277 a_189936_651879# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8278 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8279 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8280 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8281 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8282 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8283 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8284 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8285 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8286 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8287 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8288 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8289 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8290 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8291 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8292 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8293 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8294 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8295 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8296 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8297 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8298 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8299 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8300 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8301 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8302 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8303 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8304 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_434420_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8305 a_443850_641883# a_441720_645346# mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8306 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8307 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8308 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8309 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8310 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8311 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8312 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8313 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8314 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8315 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_434420_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8316 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8317 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8318 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D66 vssd1 io_analog[8] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X8319 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8320 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8321 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8322 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8323 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8324 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8325 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8326 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8327 a_203650_645683# a_201520_649146# mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8328 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8329 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8330 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8331 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8332 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8333 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8334 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8335 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8336 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8337 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8338 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8339 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8340 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8341 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8342 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8343 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8344 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8345 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8346 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8347 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8348 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8349 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8350 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8351 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8352 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8353 vccd1 io_analog[1] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X8354 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8355 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8356 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8357 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8358 vssd1 mpw5_submission_1/cmirror_channel_0/I_in_channel sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8359 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8360 mpw5_submission_1/eigth_mirror_0/I_In mpw5_submission_1/isource_0/VM22D a_171016_648702# vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8361 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8362 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8363 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8364 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8365 mpw5_submission_0/eigth_mirror_0/I_In mpw5_submission_0/isource_0/VM22D a_411216_644902# vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8366 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8367 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8368 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8369 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8370 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8371 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8372 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X8373 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8374 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8375 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_188820_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8376 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D67 io_analog[8] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X8377 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8378 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8379 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8380 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8381 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8382 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8383 a_430136_648079# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8384 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8385 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8386 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X8387 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8388 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8389 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8390 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8391 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8392 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8393 mpw5_submission_0/tia_core_0/VM31D mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8394 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8395 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8396 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8397 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8398 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8399 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8400 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8401 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8402 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8403 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8404 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8405 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8406 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8407 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8408 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8409 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8410 a_464438_656600# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8411 vssd1 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X8412 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8413 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8414 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8415 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8416 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8417 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8418 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8419 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8420 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8421 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8422 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8423 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8424 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8425 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8426 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8427 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8428 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8429 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8430 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8431 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8432 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8433 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8434 a_189446_646296# a_171016_648702# vssd1 sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X8435 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8436 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8437 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8438 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8439 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8440 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8441 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8442 io_analog[0] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X8443 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8444 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8445 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8446 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8447 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8448 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8449 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8450 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8451 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8452 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8453 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8454 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8455 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8456 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_191520_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8457 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8458 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8459 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8460 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8461 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8462 mpw5_submission_1/eigth_mirror_0/I_In mpw5_submission_1/isource_0/VM22D a_171016_648702# vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8463 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8464 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8465 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8466 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8467 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8468 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8469 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8470 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8471 a_195570_640623# mpw5_submission_1/eigth_mirror_0/I_In mpw5_submission_1/eigth_mirror_0/I_In vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8472 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8473 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X8474 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8475 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8476 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8477 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8478 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8479 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8480 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8481 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8482 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8483 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X8484 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8485 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8486 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8487 a_424970_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8488 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8489 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8490 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8491 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8492 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8493 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8494 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8495 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8496 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8497 mpw5_submission_1/tia_core_0/VM31D mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8498 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8499 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8500 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8501 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8502 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8503 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X8504 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8505 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8506 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8507 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8508 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8509 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8510 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8511 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8512 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8513 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8514 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8515 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8516 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8517 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8518 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8519 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8520 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8521 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8522 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8523 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8524 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8525 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8526 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8527 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8528 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8529 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8530 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8531 a_194220_640623# mpw5_submission_1/eigth_mirror_0/I_In mpw5_submission_1/cmirror_channel_0/I_in_channel vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8532 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8533 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8534 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8535 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8536 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8537 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8538 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8539 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8540 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8541 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8542 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8543 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8544 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8545 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8546 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8547 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8548 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8549 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_192870_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8550 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8551 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8552 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8553 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8554 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8555 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8556 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8557 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8558 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8559 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8560 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8561 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8562 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8563 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8564 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8565 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8566 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8567 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8568 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8569 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8570 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8571 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8572 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8573 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8574 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8575 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8576 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8577 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8578 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8579 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8580 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8581 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8582 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8583 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8584 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8585 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8586 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8587 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8588 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8589 a_171016_648702# mpw5_submission_1/isource_0/VM22D mpw5_submission_1/eigth_mirror_0/I_In vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8590 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8591 mpw5_submission_1/tia_core_0/VM31D mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8592 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8593 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8594 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/InputRef mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8595 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X8596 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X8597 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_194220_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8598 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8599 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8600 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8601 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8602 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8603 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8604 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8605 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8606 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8607 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8608 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8609 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8610 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8611 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8612 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8613 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8614 mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8615 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8616 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8617 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM31D mpw5_submission_0/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8618 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8619 vssd1 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM5D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8620 a_203370_649243# a_201520_649146# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8621 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8622 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8623 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8624 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8625 vccd1 io_analog[0] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X8626 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8627 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8628 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8629 mpw5_submission_1/isource_0/VM12G mpw5_submission_1/isource_0/VM14D vccd1 mpw5_submission_1/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8630 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8631 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8632 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8633 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8634 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8635 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8636 vccd1 vssd1 mpw5_submission_1/tia_core_0/Out_2 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8637 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8638 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8639 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8640 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8641 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8642 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8643 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8644 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8645 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8646 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8647 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8648 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_190170_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8649 vssd1 vccd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8650 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8651 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8652 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8653 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8654 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8655 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8656 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8657 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8658 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8659 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8660 a_441920_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8661 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8662 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8663 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8664 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8665 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8666 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8667 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8668 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8669 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8670 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8671 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8672 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8673 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8674 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8675 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8676 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8677 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8678 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8679 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8680 a_443570_645443# a_441720_645346# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8681 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8682 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8683 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8684 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8685 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8686 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8687 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8688 mpw5_submission_0/tia_core_0/VM31D mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8689 a_194220_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8690 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8691 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8692 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_191520_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8693 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8694 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8695 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8696 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8697 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8698 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8699 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8700 a_430136_645809# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8701 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8702 a_202298_647480# mpw5_submission_1/cmirror_channel_0/I_in_channel vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8703 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X8704 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D68 io_analog[2] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X8705 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM31D mpw5_submission_0/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8706 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_430370_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8707 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8708 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8709 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8710 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8711 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8712 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8713 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8714 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8715 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8716 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8717 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8718 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8719 vccd1 vssd1 mpw5_submission_0/tia_core_0/Out_2 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8720 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8721 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8722 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8723 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8724 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8725 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8726 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8727 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8728 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8729 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8730 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8731 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8732 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8733 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8734 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8735 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8736 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8737 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8738 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8739 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8740 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8741 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8742 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8743 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8744 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8745 vccd1 vssd1 mpw5_submission_1/tia_core_0/VM31D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8746 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8747 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8748 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8749 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8750 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8751 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8752 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8753 a_192870_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8754 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8755 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8756 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8757 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8758 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8759 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8760 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8761 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8762 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8763 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8764 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8765 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8766 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8767 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8768 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8769 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8770 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8771 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8772 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8773 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8774 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8775 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8776 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8777 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8778 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D69 vssd1 io_analog[8] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X8779 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8780 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8781 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8782 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8783 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8784 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8785 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8786 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8787 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8788 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8789 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8790 a_184770_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8791 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8792 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8793 mpw5_submission_0/outd_0/V_da1_P vccd1 vssd1 sky130_fd_pr__res_high_po_2p85 l=6e+06u
X8794 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8795 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8796 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8797 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8798 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8799 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8800 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8801 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8802 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8803 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8804 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8805 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8806 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8807 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8808 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8809 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8810 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8811 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8812 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8813 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8814 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8815 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8816 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8817 a_424970_636823# mpw5_submission_0/eigth_mirror_0/I_In mpw5_submission_0/eigth_mirror_0/I_out_7 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8818 mpw5_submission_1/isource_0/VM12G mpw5_submission_1/isource_0/VM14D vccd1 mpw5_submission_1/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8819 a_430136_648079# mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM14D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X8820 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8821 a_189936_651879# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8822 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8823 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8824 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8825 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8826 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8827 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8828 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8829 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8830 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8831 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8832 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8833 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8834 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8835 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8836 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8837 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8838 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8839 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8840 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8841 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8842 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8843 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8844 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8845 a_189936_660919# mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM9D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X8846 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8847 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8848 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8849 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8850 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8851 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8852 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8853 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8854 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8855 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8856 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8857 mpw5_submission_0/isource_0/VM12G mpw5_submission_0/isource_0/VM14D vccd1 mpw5_submission_0/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8858 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8859 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8860 mpw5_submission_0/eigth_mirror_0/I_out_3 mpw5_submission_0/eigth_mirror_0/I_In a_430370_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8861 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8862 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8863 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8864 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8865 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8866 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8867 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8868 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8869 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8870 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8871 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8872 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8873 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8874 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8875 mpw5_submission_0/eigth_mirror_0/I_In mpw5_submission_0/eigth_mirror_0/I_In a_435770_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8876 vccd1 mpw5_submission_1/isource_0/VM14D mpw5_submission_1/isource_0/VM12G mpw5_submission_1/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8877 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8878 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8879 vssd1 mpw5_submission_1/cmirror_channel_0/I_in_channel a_201458_647480# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8880 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8881 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8882 mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8883 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8884 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8885 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8886 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8887 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8888 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8889 mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/InputRef mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8890 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8891 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8892 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8893 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8894 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8895 a_189936_649609# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8896 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8897 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8898 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8899 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8900 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8901 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8902 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8903 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8904 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8905 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8906 vccd1 mpw5_submission_0/isource_0/VM14D mpw5_submission_0/isource_0/VM12G mpw5_submission_0/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8907 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8908 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8909 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8910 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8911 mpw5_submission_1/tia_core_0/Out_2 mpw5_submission_1/outd_0/InputSignal io_analog[6] io_analog[6] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8912 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8913 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8914 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8915 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8916 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8917 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8918 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8919 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8920 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8921 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8922 a_189936_651879# mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM14D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X8923 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8924 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8925 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8926 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8927 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8928 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8929 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8930 mpw5_submission_0/cmirror_channel_0/I_in_channel mpw5_submission_0/eigth_mirror_0/I_In a_434420_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8931 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8932 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8933 a_430136_648079# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8934 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8935 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8936 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8937 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8938 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8939 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8940 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8941 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8942 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8943 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8944 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8945 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8946 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8947 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8948 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8949 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8950 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8951 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8952 vssd1 mpw5_submission_0/cmirror_channel_0/I_in_channel a_442498_643680# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8953 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8954 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8955 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8956 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8957 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8958 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8959 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8960 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8961 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8962 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8963 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8964 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8965 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8966 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8967 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8968 vccd1 io_analog[0] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X8969 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8970 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8971 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8972 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8973 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8974 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8975 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8976 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8977 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8978 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8979 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8980 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8981 a_443570_645443# a_441720_645346# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X8982 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8983 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8984 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8985 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8986 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8987 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8988 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8989 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8990 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8991 mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8992 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8993 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8994 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8995 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8996 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8997 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8998 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8999 vccd1 io_analog[1] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X9000 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9001 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9002 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9003 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9004 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9005 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9006 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9007 a_195570_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9008 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9009 a_203650_645683# a_201520_649146# mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9010 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9011 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9012 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9013 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9014 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X9015 io_analog[5] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X9016 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9017 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9018 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9019 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9020 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D70 vssd1 io_analog[2] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X9021 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9022 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9023 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9024 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9025 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9026 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9027 io_analog[3] mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/tia_core_0/Out_2 io_analog[3] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9028 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9029 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9030 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9031 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9032 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9033 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9034 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9035 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9036 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9037 a_201458_647480# mpw5_submission_1/cmirror_channel_0/I_in_channel vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9038 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9039 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9040 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9041 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9042 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9043 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9044 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9045 mpw5_submission_1/cmirror_channel_0/I_in_channel mpw5_submission_1/cmirror_channel_0/I_in_channel a_200618_647480# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9046 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9047 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9048 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9049 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9050 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9051 vssd1 vccd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9052 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9053 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9054 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9055 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9056 vssd1 vccd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9057 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9058 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9059 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9060 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9061 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9062 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9063 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9064 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9065 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9066 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9067 a_203650_645683# a_201520_649146# mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9068 a_430706_642496# a_430176_644928# vssd1 sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X9069 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9070 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9071 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9072 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9073 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9074 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9075 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9076 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9077 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9078 a_201720_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9079 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9080 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9081 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9082 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9083 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9084 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9085 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9086 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9087 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9088 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9089 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9090 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9091 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9092 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9093 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9094 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9095 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9096 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9097 vssd1 mpw5_submission_0/cmirror_channel_0/I_in_channel a_440818_643680# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9098 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9099 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9100 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9101 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9102 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9103 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/InputRef mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9104 vssd1 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X9105 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9106 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9107 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9108 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9109 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9110 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9111 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9112 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9113 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9114 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9115 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9116 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9117 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_660919# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9118 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9119 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9120 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9121 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9122 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM6D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9123 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9124 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9125 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9126 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9127 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X9128 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9129 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9130 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X9131 a_411216_644902# mpw5_submission_0/isource_0/VM22D mpw5_submission_0/eigth_mirror_0/I_In vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9132 a_189936_660919# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9133 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9134 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9135 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9136 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9137 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9138 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9139 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9140 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9141 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9142 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9143 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9144 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9145 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9146 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9147 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9148 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9149 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9150 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9151 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9152 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9153 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9154 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9155 a_441658_643680# mpw5_submission_0/cmirror_channel_0/I_in_channel vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9156 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9157 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_187470_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9158 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9159 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9160 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9161 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9162 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9163 vccd1 io_analog[0] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X9164 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9165 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9166 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9167 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9168 mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9169 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9170 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9171 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9172 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9173 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9174 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9175 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9176 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9177 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9178 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9179 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9180 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9181 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9182 io_analog[4] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X9183 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9184 mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9185 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9186 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9187 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9188 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9189 mpw5_submission_1/isource_0/VM3D a_171016_648702# mpw5_submission_1/isource_0/VM22D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X9190 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9191 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9192 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9193 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9194 a_224238_660400# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9195 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9196 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9197 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9198 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9199 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9200 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9201 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9202 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9203 vccd1 io_analog[1] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X9204 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9205 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9206 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9207 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9208 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9209 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9210 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9211 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9212 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9213 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9214 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9215 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9216 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9217 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9218 vssd1 mpw5_submission_1/cmirror_channel_0/I_in_channel a_200618_647480# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9219 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9220 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9221 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9222 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_186120_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9223 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9224 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9225 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9226 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9227 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9228 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9229 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9230 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9231 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9232 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9233 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9234 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9235 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9236 a_191520_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9237 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9238 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9239 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9240 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9241 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9242 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9243 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9244 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9245 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_435770_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9246 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9247 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9248 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9249 io_analog[6] mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/tia_core_0/Out_2 io_analog[6] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9250 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9251 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9252 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9253 a_171016_648702# mpw5_submission_1/isource_0/VM22D mpw5_submission_1/eigth_mirror_0/I_In vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
D71 io_analog[3] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X9254 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9255 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9256 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9257 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9258 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9259 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9260 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9261 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9262 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9263 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9264 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9265 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9266 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9267 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9268 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9269 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9270 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9271 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9272 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9273 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9274 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9275 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9276 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9277 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9278 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9279 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9280 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9281 mpw5_submission_1/eigth_mirror_0/I_In mpw5_submission_1/eigth_mirror_0/I_In a_195570_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9282 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9283 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9284 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9285 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9286 mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9287 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9288 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9289 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9290 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9291 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9292 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9293 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9294 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9295 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9296 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9297 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9298 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9299 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9300 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9301 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9302 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9303 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9304 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9305 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9306 mpw5_submission_1/outd_0/V_da2_N vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X9307 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9308 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9309 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9310 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9311 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9312 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9313 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_434420_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9314 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9315 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9316 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9317 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9318 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9319 vccd1 a_441720_645346# a_441920_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9320 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9321 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9322 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9323 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9324 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9325 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9326 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9327 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9328 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9329 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9330 io_analog[4] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X9331 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9332 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9333 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9334 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9335 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9336 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9337 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9338 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9339 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9340 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9341 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9342 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9343 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9344 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9345 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9346 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9347 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9348 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9349 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9350 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9351 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9352 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9353 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9354 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9355 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9356 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9357 mpw5_submission_1/cmirror_channel_0/I_in_channel mpw5_submission_1/eigth_mirror_0/I_In a_194220_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9358 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9359 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9360 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9361 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9362 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9363 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9364 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9365 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9366 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9367 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9368 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9369 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9370 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9371 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9372 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9373 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9374 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9375 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9376 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_433070_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9377 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9378 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9379 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9380 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9381 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9382 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9383 a_189936_651879# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9384 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9385 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9386 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9387 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X9388 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X9389 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9390 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9391 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9392 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_188820_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9393 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9394 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9395 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9396 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9397 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9398 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9399 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9400 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9401 mpw5_submission_0/tia_core_0/Out_2 mpw5_submission_0/outd_0/InputSignal io_analog[3] io_analog[3] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
D72 vssd1 io_analog[7] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X9402 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9403 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9404 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9405 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9406 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9407 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9408 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9409 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9410 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D73 io_analog[8] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X9411 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9412 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9413 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9414 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9415 mpw5_submission_1/tia_core_0/VM31D mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9416 mpw5_submission_0/tia_core_0/VM5D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9417 mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/InputRef mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9418 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9419 a_224238_660400# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9420 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9421 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9422 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9423 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9424 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9425 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9426 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9427 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9428 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9429 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9430 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9431 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9432 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9433 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9434 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM31D mpw5_submission_1/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9435 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_434420_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9436 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9437 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9438 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9439 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9440 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9441 mpw5_submission_1/isource_0/VM22D a_171016_648702# mpw5_submission_1/isource_0/VM3D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X9442 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9443 mpw5_submission_0/outd_0/InputSignal io_analog[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9444 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9445 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_187470_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9446 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9447 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9448 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9449 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9450 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9451 vccd1 mpw5_submission_1/isource_0/VM14D mpw5_submission_1/isource_0/VM12G mpw5_submission_1/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9452 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9453 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9454 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9455 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9456 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9457 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9458 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9459 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9460 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9461 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9462 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9463 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9464 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9465 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9466 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9467 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9468 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9469 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9470 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9471 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9472 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9473 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9474 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9475 mpw5_submission_0/tia_core_0/VM36D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM39D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9476 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9477 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9478 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9479 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9480 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9481 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9482 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9483 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9484 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9485 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9486 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9487 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9488 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9489 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9490 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9491 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9492 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9493 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9494 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9495 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9496 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9497 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9498 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9499 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9500 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9501 a_188820_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9502 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9503 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9504 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9505 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9506 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9507 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9508 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9509 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9510 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9511 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9512 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9513 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9514 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9515 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9516 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9517 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9518 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9519 vccd1 io_analog[0] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X9520 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9521 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9522 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9523 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9524 mpw5_submission_1/eigth_mirror_0/I_In mpw5_submission_1/isource_0/VM22D a_171016_648702# vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9525 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9526 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9527 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9528 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9529 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9530 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9531 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9532 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9533 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9534 a_203370_649243# a_201520_649146# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9535 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9536 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9537 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9538 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9539 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9540 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9541 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9542 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9543 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9544 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9545 io_analog[4] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X9546 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9547 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9548 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9549 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9550 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9551 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9552 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9553 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9554 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9555 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9556 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9557 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9558 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9559 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9560 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9561 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9562 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9563 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9564 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9565 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9566 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9567 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9568 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9569 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9570 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9571 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9572 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9573 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9574 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9575 vccd1 vssd1 mpw5_submission_0/tia_core_0/VM31D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9576 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9577 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9578 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9579 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9580 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9581 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9582 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9583 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9584 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9585 a_188820_640623# mpw5_submission_1/eigth_mirror_0/I_In mpw5_submission_1/eigth_mirror_0/I_out_4 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9586 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9587 mpw5_submission_1/tia_core_0/VM31D vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9588 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9589 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9590 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9591 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9592 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9593 a_195570_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9594 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9595 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9596 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9597 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9598 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9599 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9600 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9601 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9602 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9603 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9604 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9605 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9606 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9607 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9608 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9609 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9610 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9611 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9612 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9613 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9614 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9615 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9616 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9617 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9618 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9619 vssd1 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X9620 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9621 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9622 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9623 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9624 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9625 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9626 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9627 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9628 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9629 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D74 io_analog[0] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X9630 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9631 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9632 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9633 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9634 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9635 vssd1 vccd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9636 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9637 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9638 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9639 a_424970_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9640 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9641 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9642 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9643 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9644 mpw5_submission_1/tia_core_0/Out_2 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9645 vccd1 mpw5_submission_1/isource_0/VM14D mpw5_submission_1/isource_0/VM12G mpw5_submission_1/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9646 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9647 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9648 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9649 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9650 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9651 mpw5_submission_1/outd_0/InputSignal io_analog[6] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9652 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9653 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9654 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9655 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9656 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9657 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9658 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9659 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9660 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9661 a_430136_654859# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9662 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9663 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM6D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9664 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9665 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9666 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9667 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9668 mpw5_submission_0/eigth_mirror_0/I_out_7 mpw5_submission_0/eigth_mirror_0/I_In a_424970_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9669 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9670 mpw5_submission_1/tia_core_0/VM31D mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9671 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9672 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9673 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9674 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9675 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9676 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9677 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9678 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9679 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9680 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9681 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9682 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9683 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9684 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9685 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9686 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D75 io_analog[0] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X9687 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9688 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9689 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9690 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9691 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9692 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9693 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9694 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9695 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9696 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9697 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9698 mpw5_submission_1/isource_0/VM12G mpw5_submission_1/isource_0/VM14D vccd1 mpw5_submission_1/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9699 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9700 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9701 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9702 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9703 a_431720_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9704 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9705 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9706 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9707 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9708 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9709 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9710 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9711 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9712 vccd1 io_analog[5] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X9713 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9714 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9715 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9716 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X9717 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9718 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9719 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9720 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9721 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9722 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9723 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9724 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9725 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9726 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9727 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9728 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9729 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9730 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9731 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9732 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9733 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9734 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9735 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9736 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9737 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9738 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9739 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM31D mpw5_submission_1/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9740 mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9741 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9742 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9743 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9744 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9745 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9746 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9747 a_443850_641883# a_441720_645346# mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9748 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9749 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_657119# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9750 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9751 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9752 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9753 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9754 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9755 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9756 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9757 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9758 mpw5_submission_1/tia_core_0/VM31D mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9759 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9760 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9761 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9762 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9763 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9764 a_430136_657119# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9765 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9766 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9767 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9768 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9769 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9770 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9771 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9772 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9773 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9774 a_203370_649243# a_201520_649146# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9775 a_430706_642496# a_431236_644928# vssd1 sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X9776 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9777 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9778 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9779 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9780 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9781 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9782 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9783 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9784 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9785 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9786 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9787 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9788 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9789 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9790 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9791 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9792 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9793 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9794 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9795 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9796 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9797 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9798 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9799 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9800 mpw5_submission_0/isource_0/VM22D a_411216_644902# mpw5_submission_0/isource_0/VM3D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X9801 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9802 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9803 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9804 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9805 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9806 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9807 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9808 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9809 a_189936_651879# mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM14D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X9810 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9811 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9812 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9813 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9814 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9815 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9816 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9817 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9818 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9819 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9820 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9821 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9822 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X9823 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9824 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9825 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9826 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9827 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9828 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9829 a_203370_649243# a_201520_649146# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9830 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9831 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9832 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X9833 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9834 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9835 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9836 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9837 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9838 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9839 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9840 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9841 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9842 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9843 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9844 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9845 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9846 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9847 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9848 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9849 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X9850 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9851 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9852 mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9853 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9854 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9855 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9856 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9857 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9858 vssd1 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X9859 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9860 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9861 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9862 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9863 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9864 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9865 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9866 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9867 mpw5_submission_0/tia_core_0/VM31D mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9868 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9869 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9870 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9871 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9872 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9873 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9874 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9875 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D76 vssd1 io_analog[1] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X9876 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9877 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9878 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9879 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9880 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9881 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9882 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9883 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9884 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9885 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9886 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9887 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9888 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9889 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9890 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9891 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9892 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9893 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9894 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9895 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9896 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9897 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9898 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9899 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9900 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9901 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9902 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9903 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9904 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9905 vccd1 io_analog[5] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X9906 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9907 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9908 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9909 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9910 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9911 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9912 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9913 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9914 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9915 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9916 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9917 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9918 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9919 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9920 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9921 mpw5_submission_0/outd_0/InputSignal io_analog[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9922 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9923 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9924 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9925 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9926 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9927 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9928 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9929 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9930 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9931 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9932 a_430136_648079# mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM14D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
D77 io_analog[8] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X9933 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9934 a_189936_651879# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9935 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9936 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9937 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9938 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9939 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X9940 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9941 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9942 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X9943 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9944 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9945 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9946 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9947 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9948 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9949 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9950 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9951 a_434420_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9952 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9953 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9954 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9955 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9956 mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9957 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9958 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9959 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9960 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9961 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9962 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X9963 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9964 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9965 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9966 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9967 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9968 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9969 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9970 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9971 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9972 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9973 a_427116_648806# a_427646_651238# vssd1 sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X9974 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9975 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9976 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9977 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9978 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9979 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9980 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9981 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9982 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9983 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9984 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9985 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9986 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9987 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9988 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9989 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9990 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9991 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9992 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9993 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9994 vccd1 io_analog[7] mpw5_submission_0/tia_core_0/Disable_TIA_B vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=1e+06u
X9995 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9996 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9997 io_analog[1] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X9998 vssd1 vccd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9999 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10000 mpw5_submission_0/tia_core_0/VM6D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10001 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10002 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10003 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10004 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10005 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10006 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10007 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10008 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10009 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10010 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10011 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10012 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10013 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10014 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10015 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10016 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10017 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10018 io_analog[4] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X10019 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10020 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10021 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10022 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10023 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10024 vccd1 vssd1 mpw5_submission_0/tia_core_0/Out_2 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10025 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10026 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10027 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10028 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_188820_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10029 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10030 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10031 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10032 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10033 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10034 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10035 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10036 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10037 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10038 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10039 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10040 a_430136_648079# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10041 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10042 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10043 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10044 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10045 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X10046 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X10047 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10048 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10049 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10050 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10051 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10052 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10053 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10054 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10055 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10056 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10057 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10058 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X10059 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10060 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10061 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10062 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10063 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X10064 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10065 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10066 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10067 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10068 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10069 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10070 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10071 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10072 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10073 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10074 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10075 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10076 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10077 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10078 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10079 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10080 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10081 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10082 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10083 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10084 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10085 vssd1 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X10086 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10087 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10088 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10089 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10090 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10091 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10092 a_203370_649243# a_201520_649146# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10093 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10094 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10095 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10096 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10097 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10098 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10099 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10100 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10101 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10102 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10103 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10104 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10105 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10106 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10107 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10108 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10109 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10110 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10111 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10112 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10113 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10114 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10115 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10116 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10117 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10118 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10119 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10120 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10121 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10122 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10123 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10124 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10125 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10126 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10127 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10128 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10129 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10130 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10131 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10132 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10133 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10134 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_424970_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10135 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10136 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10137 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10138 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10139 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10140 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10141 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10142 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10143 mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10144 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10145 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10146 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10147 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10148 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_424970_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10149 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10150 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10151 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10152 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10153 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10154 vssd1 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 sky130_fd_pr__cap_mim_m3_1 l=1.2e+07u w=1.5e+07u
X10155 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10156 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10157 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10158 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10159 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10160 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10161 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10162 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10163 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10164 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10165 a_190170_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10166 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10167 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10168 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10169 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10170 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10171 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_660919# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10172 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10173 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10174 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10175 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10176 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10177 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10178 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10179 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10180 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10181 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10182 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10183 vccd1 io_analog[4] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X10184 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10185 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10186 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10187 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10188 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10189 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10190 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10191 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10192 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10193 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10194 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10195 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10196 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10197 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10198 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10199 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10200 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10201 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_426320_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10202 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10203 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10204 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10205 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10206 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10207 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10208 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10209 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10210 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10211 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10212 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10213 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10214 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10215 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10216 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10217 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10218 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10219 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10220 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10221 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10222 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10223 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10224 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10225 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10226 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10227 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10228 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10229 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10230 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10231 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10232 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10233 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10234 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D78 vssd1 io_analog[0] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X10235 mpw5_submission_1/tia_core_0/VM6D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10236 vssd1 mpw5_submission_0/isource_0/VM3G mpw5_submission_0/isource_0/VM3D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X10237 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10238 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10239 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10240 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10241 vssd1 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM36D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10242 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10243 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM36D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10244 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10245 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10246 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10247 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10248 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10249 a_191520_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10250 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10251 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10252 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10253 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10254 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10255 a_435770_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10256 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10257 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10258 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10259 vccd1 mpw5_submission_1/outd_0/V_da2_P vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X10260 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10261 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10262 mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10263 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10264 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10265 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10266 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10267 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10268 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10269 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10270 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10271 a_189936_649609# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10272 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10273 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10274 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10275 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10276 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10277 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10278 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10279 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10280 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10281 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10282 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10283 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10284 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10285 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10286 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10287 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10288 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10289 mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10290 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10291 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10292 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10293 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10294 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10295 io_analog[0] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X10296 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10297 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10298 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10299 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10300 a_171016_648702# mpw5_submission_1/isource_0/VM22D mpw5_submission_1/eigth_mirror_0/I_In vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10301 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10302 vccd1 a_201520_649146# a_201720_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10303 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X10304 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10305 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10306 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10307 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10308 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10309 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10310 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10311 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10312 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10313 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10314 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10315 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10316 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10317 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10318 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10319 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10320 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10321 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10322 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10323 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10324 vccd1 a_441720_645346# a_441920_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10325 vccd1 vssd1 mpw5_submission_1/tia_core_0/Out_2 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10326 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10327 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10328 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10329 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10330 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10331 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10332 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10333 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10334 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10335 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10336 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10337 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10338 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10339 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10340 a_190170_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10341 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10342 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10343 mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10344 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10345 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10346 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10347 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10348 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10349 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10350 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10351 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10352 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10353 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10354 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10355 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10356 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10357 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10358 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10359 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10360 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10361 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10362 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM36D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10363 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10364 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_645809# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10365 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10366 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10367 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10368 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10369 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10370 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10371 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10372 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10373 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_191520_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10374 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10375 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10376 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10377 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10378 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10379 a_430136_645809# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10380 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10381 a_200618_647480# mpw5_submission_1/cmirror_channel_0/I_in_channel vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10382 a_184770_640623# mpw5_submission_1/eigth_mirror_0/I_In mpw5_submission_1/eigth_mirror_0/I_out_7 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10383 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10384 mpw5_submission_1/tia_core_0/VM5D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10385 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10386 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10387 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10388 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10389 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10390 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10391 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10392 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10393 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10394 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10395 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10396 mpw5_submission_0/outd_0/InputSignal io_analog[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10397 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10398 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10399 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10400 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10401 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10402 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10403 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10404 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10405 a_443570_645443# a_441720_645346# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10406 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10407 mpw5_submission_1/isource_0/VM12G mpw5_submission_1/isource_0/VM14D vccd1 mpw5_submission_1/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10408 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10409 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10410 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10411 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10412 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10413 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10414 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10415 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10416 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X10417 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10418 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10419 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10420 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10421 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10422 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10423 mpw5_submission_0/tia_core_0/VM6D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10424 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10425 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10426 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10427 mpw5_submission_1/eigth_mirror_0/I_In mpw5_submission_1/eigth_mirror_0/I_In a_195570_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10428 mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10429 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10430 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10431 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10432 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10433 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10434 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10435 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10436 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10437 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10438 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10439 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10440 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10441 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10442 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10443 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10444 mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10445 vssd1 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 sky130_fd_pr__cap_mim_m3_1 l=1.2e+07u w=1.5e+07u
X10446 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10447 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10448 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10449 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10450 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10451 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10452 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10453 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10454 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10455 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10456 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10457 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10458 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10459 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10460 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10461 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10462 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10463 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10464 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10465 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10466 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10467 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10468 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10469 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10470 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D79 io_analog[7] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X10471 mpw5_submission_0/outd_0/V_da2_P vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X10472 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10473 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10474 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10475 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10476 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10477 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10478 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10479 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10480 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10481 mpw5_submission_1/cmirror_channel_0/I_in_channel mpw5_submission_1/eigth_mirror_0/I_In a_194220_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10482 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10483 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10484 a_189936_651879# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10485 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10486 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10487 a_203650_645683# a_201520_649146# mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10488 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10489 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10490 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10491 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10492 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10493 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10494 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10495 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10496 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10497 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10498 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10499 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10500 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10501 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10502 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10503 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10504 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10505 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10506 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10507 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10508 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10509 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10510 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10511 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10512 a_203370_649243# a_201520_649146# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10513 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10514 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10515 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10516 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10517 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10518 a_201458_647480# mpw5_submission_1/cmirror_channel_0/I_in_channel vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10519 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10520 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10521 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10522 vccd1 io_analog[4] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X10523 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10524 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10525 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10526 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10527 mpw5_submission_1/tia_core_0/VM31D mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10528 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10529 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10530 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10531 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10532 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10533 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10534 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_649609# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10535 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10536 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D80 io_analog[3] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X10537 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10538 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10539 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10540 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10541 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10542 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10543 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10544 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10545 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10546 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10547 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10548 vccd1 io_analog[1] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X10549 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10550 a_189936_649609# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10551 mpw5_submission_0/outd_0/InputSignal io_analog[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10552 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10553 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10554 a_195570_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10555 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10556 vccd1 io_analog[5] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X10557 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10558 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10559 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10560 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10561 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10562 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10563 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10564 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10565 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10566 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10567 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10568 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10569 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10570 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10571 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10572 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10573 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10574 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10575 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10576 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10577 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10578 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10579 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10580 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10581 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10582 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10583 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10584 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10585 mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10586 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10587 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10588 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10589 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10590 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10591 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10592 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10593 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10594 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10595 mpw5_submission_1/outd_0/InputSignal io_analog[6] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10596 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10597 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10598 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10599 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10600 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10601 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D81 vssd1 io_analog[7] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X10602 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10603 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10604 a_194220_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10605 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10606 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10607 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10608 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10609 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10610 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10611 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10612 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10613 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10614 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10615 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10616 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10617 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10618 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10619 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10620 a_190506_646296# a_189976_648728# vssd1 sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X10621 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10622 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10623 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10624 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10625 mpw5_submission_0/outd_0/V_da1_P vccd1 vssd1 sky130_fd_pr__res_high_po_2p85 l=6e+06u
X10626 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10627 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10628 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10629 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10630 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10631 a_428176_648806# a_427646_651238# vssd1 sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X10632 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10633 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10634 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10635 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10636 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D82 vssd1 io_analog[0] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X10637 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10638 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10639 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10640 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10641 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10642 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10643 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10644 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10645 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM31D mpw5_submission_0/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10646 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10647 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10648 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10649 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10650 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10651 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10652 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10653 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10654 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_195570_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10655 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10656 a_192870_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10657 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10658 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10659 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D83 vssd1 io_analog[1] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X10660 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10661 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10662 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10663 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10664 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10665 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10666 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10667 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10668 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10669 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10670 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10671 a_185856_652606# a_185326_655038# vssd1 sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X10672 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10673 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10674 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10675 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10676 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10677 a_431720_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10678 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10679 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10680 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10681 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10682 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10683 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10684 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10685 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10686 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10687 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10688 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X10689 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10690 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10691 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10692 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10693 vssd1 mpw5_submission_1/cmirror_channel_0/I_in_channel a_200618_647480# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10694 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10695 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10696 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10697 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10698 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10699 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10700 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10701 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10702 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10703 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10704 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10705 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10706 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10707 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10708 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_429020_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10709 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10710 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10711 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10712 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10713 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10714 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10715 vccd1 io_analog[4] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X10716 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10717 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10718 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10719 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10720 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10721 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10722 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10723 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10724 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10725 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10726 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10727 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10728 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10729 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10730 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10731 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10732 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D84 vssd1 io_analog[0] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X10733 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10734 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10735 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10736 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10737 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10738 vccd1 io_analog[5] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X10739 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10740 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10741 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10742 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10743 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10744 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10745 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10746 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10747 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10748 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10749 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10750 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10751 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10752 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10753 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10754 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10755 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10756 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10757 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10758 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10759 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10760 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10761 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10762 mpw5_submission_0/eigth_mirror_0/I_out_7 mpw5_submission_0/eigth_mirror_0/I_In a_424970_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10763 mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/InputRef mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10764 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10765 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10766 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10767 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10768 vssd1 vccd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10769 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10770 vccd1 mpw5_submission_0/outd_0/V_da2_P vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X10771 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10772 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10773 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10774 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10775 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10776 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10777 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10778 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10779 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10780 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10781 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10782 vccd1 mpw5_submission_0/isource_0/VM14D mpw5_submission_0/isource_0/VM12G mpw5_submission_0/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10783 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10784 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10785 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10786 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10787 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10788 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10789 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10790 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10791 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10792 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10793 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10794 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10795 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10796 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10797 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10798 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10799 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10800 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10801 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10802 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10803 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10804 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10805 mpw5_submission_0/tia_core_0/VM31D vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10806 vccd1 mpw5_submission_1/outd_0/V_da2_N vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X10807 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10808 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10809 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10810 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10811 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10812 mpw5_submission_1/tia_core_0/VM36D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM39D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10813 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10814 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10815 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10816 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10817 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10818 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10819 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10820 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10821 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10822 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10823 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10824 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10825 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10826 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10827 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10828 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10829 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10830 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10831 io_analog[1] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X10832 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10833 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM31D mpw5_submission_1/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10834 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10835 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10836 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10837 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10838 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10839 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10840 a_186120_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10841 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10842 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10843 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10844 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10845 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10846 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10847 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10848 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10849 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10850 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10851 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10852 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10853 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10854 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10855 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10856 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X10857 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10858 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10859 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10860 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10861 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10862 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10863 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10864 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10865 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10866 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10867 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10868 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10869 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10870 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10871 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10872 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10873 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10874 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10875 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10876 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10877 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10878 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10879 vccd1 vssd1 mpw5_submission_1/tia_core_0/Out_2 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10880 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10881 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10882 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10883 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10884 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10885 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10886 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10887 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10888 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10889 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10890 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10891 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10892 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10893 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10894 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10895 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10896 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10897 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10898 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10899 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10900 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10901 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10902 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10903 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10904 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10905 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10906 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10907 a_195570_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10908 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10909 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10910 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10911 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10912 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10913 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10914 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10915 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10916 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10917 a_202298_647480# mpw5_submission_1/cmirror_channel_0/I_in_channel mpw5_submission_1/cmirror_channel_0/TIA_I_Bias2 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
R3 vccd1 io_clamp_high[0] sky130_fd_pr__res_generic_m3 w=1.1e+07u l=250000u
X10918 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10919 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10920 a_434420_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10921 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10922 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10923 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10924 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10925 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10926 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10927 mpw5_submission_0/outd_0/InputSignal io_analog[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10928 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10929 a_192870_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10930 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10931 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10932 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10933 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10934 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10935 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10936 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10937 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10938 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10939 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10940 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10941 vccd1 a_441720_645346# a_441920_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10942 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10943 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10944 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10945 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10946 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10947 a_430136_648079# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10948 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10949 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10950 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10951 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10952 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10953 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10954 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10955 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10956 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10957 mpw5_submission_0/tia_core_0/VM31D mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10958 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10959 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10960 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10961 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10962 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10963 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10964 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10965 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10966 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10967 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10968 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10969 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10970 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10971 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10972 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10973 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10974 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10975 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10976 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10977 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X10978 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10979 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10980 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10981 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10982 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10983 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10984 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10985 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10986 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10987 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10988 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10989 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10990 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10991 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10992 io_analog[3] mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM5D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10993 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10994 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10995 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10996 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM6D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10997 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10998 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10999 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_188820_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11000 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11001 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11002 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11003 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11004 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11005 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11006 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11007 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11008 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11009 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11010 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11011 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11012 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11013 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11014 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11015 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X11016 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11017 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11018 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11019 vccd1 io_analog[4] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X11020 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11021 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11022 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11023 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11024 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11025 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11026 mpw5_submission_0/tia_core_0/VM5D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11027 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11028 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11029 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11030 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D85 vssd1 io_analog[2] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X11031 mpw5_submission_0/outd_0/V_da2_N vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X11032 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11033 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11034 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11035 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11036 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11037 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11038 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11039 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11040 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11041 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11042 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11043 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11044 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11045 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11046 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11047 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias2 mpw5_submission_0/cmirror_channel_0/I_in_channel a_442498_643680# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11048 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11049 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11050 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11051 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11052 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11053 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_187470_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11054 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11055 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11056 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11057 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11058 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11059 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11060 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11061 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11062 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11063 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11064 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11065 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11066 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11067 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11068 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11069 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11070 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11071 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11072 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11073 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11074 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11075 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11076 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11077 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11078 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11079 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11080 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11081 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11082 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11083 a_189936_651879# mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM14D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X11084 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11085 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X11086 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11087 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11088 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11089 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11090 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11091 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11092 mpw5_submission_1/isource_0/VM22D a_171016_648702# mpw5_submission_1/isource_0/VM3D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X11093 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11094 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11095 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11096 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11097 mpw5_submission_1/outd_0/V_da1_N vccd1 vssd1 sky130_fd_pr__res_high_po_2p85 l=6e+06u
X11098 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11099 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11100 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11101 mpw5_submission_0/isource_0/VM22D a_411216_644902# mpw5_submission_0/isource_0/VM3D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X11102 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11103 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11104 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11105 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11106 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11107 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11108 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11109 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11110 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11111 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11112 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11113 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11114 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_186120_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11115 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11116 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11117 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11118 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11119 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11120 a_443850_641883# a_441720_645346# mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11121 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11122 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11123 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11124 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11125 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11126 mpw5_submission_0/tia_core_0/VM36D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM39D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11127 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11128 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11129 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11130 vssd1 vccd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X11131 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11132 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11133 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11134 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11135 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11136 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11137 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11138 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_424970_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11139 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11140 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11141 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11142 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11143 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11144 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11145 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11146 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11147 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11148 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11149 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11150 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11151 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11152 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11153 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11154 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11155 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11156 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11157 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11158 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11159 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11160 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11161 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11162 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11163 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11164 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11165 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11166 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11167 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11168 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11169 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11170 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11171 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11172 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X11173 a_189936_658659# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X11174 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11175 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11176 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11177 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11178 mpw5_submission_1/eigth_mirror_0/I_out_7 mpw5_submission_1/eigth_mirror_0/I_In a_184770_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11179 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11180 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11181 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11182 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11183 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11184 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11185 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11186 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11187 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11188 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11189 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11190 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11191 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_426320_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11192 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11193 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11194 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11195 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11196 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11197 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11198 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11199 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11200 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11201 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11202 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11203 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11204 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11205 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11206 vssd1 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM6D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11207 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11208 a_203370_649243# a_201520_649146# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11209 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11210 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11211 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11212 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11213 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11214 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11215 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11216 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11217 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11218 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11219 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11220 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11221 vssd1 mpw5_submission_0/cmirror_channel_0/I_in_channel a_442498_643680# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11222 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11223 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11224 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11225 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11226 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11227 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11228 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11229 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11230 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11231 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11232 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11233 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11234 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11235 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11236 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11237 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11238 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11239 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11240 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11241 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11242 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11243 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11244 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11245 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11246 vccd1 io_analog[1] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X11247 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_424970_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11248 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11249 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11250 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11251 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D86 io_analog[0] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X11252 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11253 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11254 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11255 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11256 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11257 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11258 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11259 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11260 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11261 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11262 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11263 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11264 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11265 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11266 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_654859# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X11267 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11268 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11269 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11270 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11271 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11272 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11273 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11274 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11275 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11276 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11277 a_430136_654859# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X11278 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11279 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11280 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11281 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11282 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11283 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11284 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11285 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11286 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11287 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11288 a_190506_646296# a_191036_648728# vssd1 sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X11289 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11290 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11291 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11292 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11293 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11294 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11295 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11296 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D87 io_analog[1] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X11297 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11298 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11299 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11300 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D88 io_analog[0] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X11301 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11302 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11303 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11304 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11305 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11306 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11307 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11308 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11309 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11310 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11311 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11312 a_190170_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11313 vssd1 vccd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X11314 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11315 mpw5_submission_0/tia_core_0/VM36D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM39D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11316 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11317 mpw5_submission_0/isource_0/VM3D a_411216_644902# mpw5_submission_0/isource_0/VM22D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X11318 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11319 mpw5_submission_0/isource_0/VM3D a_411216_644902# mpw5_submission_0/isource_0/VM22D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X11320 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11321 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11322 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11323 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11324 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11325 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11326 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11327 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11328 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11329 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11330 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11331 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11332 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11333 mpw5_submission_0/eigth_mirror_0/I_out_6 mpw5_submission_0/eigth_mirror_0/I_In a_426320_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11334 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11335 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11336 a_185856_652606# a_186386_655038# vssd1 sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X11337 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11338 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11339 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11340 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11341 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11342 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D89 vssd1 io_analog[7] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X11343 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11344 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11345 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11346 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11347 a_430136_654859# mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM8D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X11348 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11349 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11350 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11351 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11352 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11353 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11354 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11355 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11356 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11357 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X11358 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11359 a_435770_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11360 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11361 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11362 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11363 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11364 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
R4 vccd1 io_clamp_high[1] sky130_fd_pr__res_generic_m3 w=1.1e+07u l=250000u
X11365 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11366 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11367 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11368 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11369 a_188820_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11370 a_430370_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11371 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11372 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11373 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11374 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11375 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11376 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11377 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11378 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11379 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_657119# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X11380 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11381 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11382 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X11383 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11384 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X11385 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11386 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11387 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11388 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11389 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11390 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11391 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11392 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11393 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11394 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11395 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11396 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11397 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11398 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11399 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11400 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11401 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11402 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11403 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11404 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11405 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11406 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11407 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11408 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11409 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11410 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11411 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11412 mpw5_submission_0/isource_0/VM12G a_424386_651238# vssd1 sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X11413 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11414 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11415 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11416 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11417 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11418 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11419 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11420 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11421 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11422 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11423 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11424 a_443850_641883# a_441720_645346# mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11425 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11426 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11427 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11428 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11429 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11430 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11431 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11432 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11433 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11434 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11435 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11436 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11437 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11438 vssd1 mpw5_submission_1/cmirror_channel_0/I_in_channel a_202298_647480# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11439 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11440 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11441 a_184770_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11442 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D90 io_analog[0] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X11443 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11444 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11445 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11446 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11447 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11448 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11449 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11450 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11451 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11452 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11453 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11454 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11455 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11456 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11457 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11458 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11459 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11460 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11461 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11462 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11463 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11464 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11465 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11466 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11467 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11468 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11469 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11470 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11471 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11472 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11473 vccd1 mpw5_submission_0/outd_0/V_da2_P vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X11474 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11475 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11476 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11477 mpw5_submission_1/outd_0/InputSignal io_analog[6] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11478 mpw5_submission_0/outd_0/V_da1_N vccd1 vssd1 sky130_fd_pr__res_high_po_2p85 l=6e+06u
X11479 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11480 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11481 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11482 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11483 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11484 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11485 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11486 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11487 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11488 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11489 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11490 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11491 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11492 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11493 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X11494 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11495 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11496 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11497 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11498 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11499 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11500 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM6D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11501 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11502 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11503 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11504 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM6D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11505 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11506 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11507 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D91 io_analog[0] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X11508 vccd1 io_analog[1] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X11509 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11510 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11511 mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11512 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11513 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11514 mpw5_submission_0/outd_0/InputSignal io_analog[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11515 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11516 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11517 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11518 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11519 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11520 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11521 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11522 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X11523 io_analog[5] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X11524 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11525 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11526 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11527 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11528 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11529 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11530 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11531 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11532 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11533 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11534 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11535 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11536 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11537 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11538 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11539 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11540 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11541 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11542 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11543 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11544 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11545 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11546 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11547 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11548 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11549 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11550 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11551 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X11552 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11553 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11554 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11555 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11556 vccd1 mpw5_submission_1/tia_core_0/Disable_TIA mpw5_submission_1/tia_core_0/Disable_TIA_B vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=1e+06u
X11557 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11558 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11559 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11560 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11561 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11562 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11563 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11564 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11565 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11566 a_189936_651879# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X11567 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11568 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11569 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11570 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11571 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11572 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11573 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11574 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11575 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11576 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11577 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11578 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11579 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11580 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11581 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11582 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11583 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11584 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11585 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11586 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X11587 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X11588 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11589 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11590 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11591 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11592 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11593 mpw5_submission_0/outd_0/V_da1_N vccd1 vssd1 sky130_fd_pr__res_high_po_2p85 l=6e+06u
X11594 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11595 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11596 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11597 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11598 a_203650_645683# a_201520_649146# mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11599 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11600 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11601 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11602 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM36D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11603 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11604 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11605 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11606 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11607 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X11608 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11609 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11610 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11611 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11612 mpw5_submission_1/outd_0/InputSignal io_analog[6] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11613 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11614 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11615 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11616 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11617 a_433070_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11618 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11619 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X11620 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11621 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11622 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11623 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11624 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11625 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X11626 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11627 a_435770_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11628 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11629 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11630 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11631 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11632 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11633 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11634 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11635 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11636 mpw5_submission_1/outd_0/InputSignal io_analog[6] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11637 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11638 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11639 a_188820_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11640 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11641 io_analog[5] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X11642 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11643 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11644 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11645 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11646 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11647 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11648 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11649 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11650 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11651 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11652 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11653 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11654 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11655 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11656 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11657 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11658 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X11659 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11660 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11661 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11662 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11663 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11664 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11665 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11666 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11667 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11668 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11669 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11670 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11671 vccd1 vssd1 mpw5_submission_0/tia_core_0/Out_2 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11672 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11673 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11674 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11675 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D92 io_analog[2] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X11676 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11677 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11678 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11679 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11680 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11681 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11682 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11683 mpw5_submission_1/tia_core_0/Out_2 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11684 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11685 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11686 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11687 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11688 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11689 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11690 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11691 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11692 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11693 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11694 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11695 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11696 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11697 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11698 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11699 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11700 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11701 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11702 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11703 a_187470_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11704 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11705 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11706 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11707 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11708 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11709 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11710 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11711 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11712 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11713 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11714 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11715 vccd1 io_analog[0] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X11716 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11717 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11718 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11719 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11720 mpw5_submission_1/outd_0/InputSignal io_analog[6] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11721 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11722 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11723 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11724 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11725 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11726 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X11727 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11728 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11729 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X11730 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11731 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11732 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11733 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11734 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11735 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11736 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11737 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11738 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11739 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11740 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11741 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11742 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11743 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11744 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11745 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11746 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11747 vssd1 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X11748 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11749 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11750 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11751 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11752 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11753 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11754 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11755 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11756 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11757 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11758 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11759 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11760 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11761 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11762 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11763 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11764 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_190170_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11765 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11766 io_analog[3] mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/tia_core_0/Out_2 io_analog[3] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11767 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11768 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11769 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11770 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11771 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11772 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11773 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11774 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11775 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11776 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11777 vccd1 io_analog[0] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X11778 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11779 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11780 mpw5_submission_1/tia_core_0/VM31D vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11781 mpw5_submission_1/tia_core_0/VM6D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11782 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11783 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11784 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11785 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11786 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11787 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11788 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11789 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11790 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11791 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11792 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11793 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11794 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11795 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11796 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11797 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11798 io_analog[4] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X11799 vccd1 mpw5_submission_0/isource_0/VM11D a_422158_661070# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X11800 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11801 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11802 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11803 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11804 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11805 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11806 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_429020_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
D93 vssd1 io_analog[7] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X11807 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11808 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11809 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11810 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11811 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11812 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11813 io_analog[0] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X11814 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11815 a_443570_645443# a_441720_645346# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11816 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11817 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11818 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11819 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11820 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11821 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11822 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11823 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11824 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11825 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11826 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11827 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11828 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11829 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11830 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11831 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11832 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X11833 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11834 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11835 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11836 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11837 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11838 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11839 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11840 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11841 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11842 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11843 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11844 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X11845 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11846 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11847 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11848 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11849 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11850 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11851 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11852 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11853 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11854 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11855 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11856 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11857 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11858 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11859 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11860 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11861 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11862 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11863 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11864 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11865 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11866 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11867 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11868 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11869 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11870 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11871 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11872 mpw5_submission_1/outd_0/V_da2_P vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X11873 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11874 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11875 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_649609# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X11876 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11877 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11878 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11879 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11880 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11881 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11882 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11883 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11884 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11885 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11886 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11887 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X11888 a_189936_649609# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X11889 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11890 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11891 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11892 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11893 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11894 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11895 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11896 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11897 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11898 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11899 mpw5_submission_0/outd_0/InputSignal io_analog[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11900 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11901 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11902 a_203370_649243# a_201520_649146# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11903 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11904 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11905 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11906 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11907 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11908 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11909 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11910 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11911 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11912 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11913 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11914 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11915 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11916 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11917 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11918 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11919 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11920 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11921 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11922 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11923 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11924 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11925 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11926 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11927 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11928 vccd1 a_201520_649146# a_201720_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11929 a_192870_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11930 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11931 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11932 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11933 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11934 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11935 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11936 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11937 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11938 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11939 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11940 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11941 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11942 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11943 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11944 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11945 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11946 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11947 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11948 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X11949 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X11950 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11951 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11952 vccd1 a_441720_645346# a_441920_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11953 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11954 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11955 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11956 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11957 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11958 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11959 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11960 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11961 a_433070_636823# mpw5_submission_0/eigth_mirror_0/I_In io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11962 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11963 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11964 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11965 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11966 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11967 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11968 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11969 a_203370_649243# a_201520_649146# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11970 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11971 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11972 mpw5_submission_1/tia_core_0/VM36D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11973 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X11974 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D94 vssd1 io_analog[1] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X11975 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11976 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11977 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11978 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11979 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11980 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11981 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11982 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11983 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11984 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11985 mpw5_submission_0/tia_core_0/VM5D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 io_analog[3] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11986 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11987 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11988 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11989 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11990 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11991 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11992 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11993 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11994 io_analog[3] mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/tia_core_0/Out_2 io_analog[3] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11995 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_645809# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X11996 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11997 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11998 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11999 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12000 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12001 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12002 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12003 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D95 io_analog[7] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X12004 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12005 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12006 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12007 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12008 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12009 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12010 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12011 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12012 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12013 mpw5_submission_1/outd_0/V_da1_P vccd1 vssd1 sky130_fd_pr__res_high_po_2p85 l=6e+06u
X12014 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12015 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12016 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12017 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12018 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12019 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12020 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12021 mpw5_submission_1/tia_core_0/VM5D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12022 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12023 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12024 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12025 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12026 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12027 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12028 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12029 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12030 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12031 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12032 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12033 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12034 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12035 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12036 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12037 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12038 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12039 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12040 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12041 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12042 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12043 a_190170_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12044 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12045 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12046 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12047 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12048 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12049 a_430136_648079# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X12050 a_422158_661070# mpw5_submission_0/isource_0/VM11D vssd1 vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X12051 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12052 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12053 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12054 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12055 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12056 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12057 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12058 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12059 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12060 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12061 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12062 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12063 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12064 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12065 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12066 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12067 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12068 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12069 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12070 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12071 a_426320_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12072 mpw5_submission_0/outd_0/InputSignal io_analog[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12073 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12074 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12075 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12076 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12077 a_443570_645443# a_441720_645346# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12078 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12079 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12080 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12081 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12082 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12083 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12084 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12085 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12086 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12087 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12088 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12089 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12090 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12091 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12092 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12093 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12094 a_190170_640623# mpw5_submission_1/eigth_mirror_0/I_In mpw5_submission_1/eigth_mirror_0/I_out_3 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12095 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12096 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12097 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM36D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12098 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12099 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12100 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12101 vccd1 vssd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X12102 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12103 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12104 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12105 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12106 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12107 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12108 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12109 mpw5_submission_0/isource_0/VM3D a_411216_644902# mpw5_submission_0/isource_0/VM22D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X12110 mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X12111 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12112 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12113 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12114 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12115 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12116 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12117 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12118 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12119 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12120 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12121 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12122 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12123 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12124 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12125 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12126 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12127 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12128 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X12129 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12130 a_424970_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12131 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12132 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12133 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12134 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12135 a_443570_645443# a_441720_645346# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12136 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12137 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12138 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12139 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12140 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12141 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12142 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12143 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12144 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12145 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12146 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12147 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12148 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12149 a_427670_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12150 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12151 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12152 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12153 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12154 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12155 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12156 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12157 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D96 vssd1 io_analog[3] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X12158 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12159 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12160 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12161 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12162 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12163 a_203650_645683# a_201520_649146# mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12164 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12165 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12166 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12167 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12168 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12169 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12170 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12171 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12172 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12173 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12174 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12175 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12176 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12177 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12178 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12179 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12180 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12181 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12182 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12183 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12184 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12185 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12186 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12187 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12188 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12189 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12190 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12191 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12192 a_443850_641883# a_441720_645346# mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12193 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12194 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12195 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12196 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12197 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12198 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12199 io_analog[6] mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/tia_core_0/Out_2 io_analog[6] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12200 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12201 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12202 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12203 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12204 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12205 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12206 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12207 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12208 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12209 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12210 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12211 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12212 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12213 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12214 a_203370_649243# a_201520_649146# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12215 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12216 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12217 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12218 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X12219 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12220 mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X12221 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12222 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12223 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12224 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12225 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12226 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12227 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12228 vssd1 vccd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X12229 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12230 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12231 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12232 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12233 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12234 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
D97 io_analog[8] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X12235 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12236 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12237 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12238 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12239 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12240 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12241 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12242 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12243 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12244 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12245 a_443850_641883# a_441720_645346# mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12246 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12247 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12248 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12249 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12250 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12251 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12252 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12253 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12254 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12255 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12256 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12257 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12258 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12259 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12260 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12261 a_431720_636823# mpw5_submission_0/eigth_mirror_0/I_In mpw5_submission_0/eigth_mirror_0/I_out_2 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12262 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12263 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12264 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12265 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12266 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224238_660400# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12267 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12268 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12269 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12270 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12271 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12272 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12273 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12274 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12275 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12276 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12277 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12278 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12279 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12280 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12281 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12282 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_654859# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X12283 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12284 mpw5_submission_0/outd_0/V_da2_N vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X12285 mpw5_submission_0/tia_core_0/VM6D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12286 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12287 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12288 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12289 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12290 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12291 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12292 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12293 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12294 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12295 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12296 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12297 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12298 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12299 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X12300 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_195570_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12301 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12302 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12303 a_441920_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12304 mpw5_submission_1/eigth_mirror_0/I_out_7 mpw5_submission_1/eigth_mirror_0/I_In a_184770_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12305 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12306 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12307 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12308 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12309 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12310 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12311 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12312 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12313 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12314 mpw5_submission_0/eigth_mirror_0/I_In mpw5_submission_0/isource_0/VM22D a_411216_644902# vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X12315 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12316 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12317 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12318 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12319 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12320 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12321 mpw5_submission_0/tia_core_0/Out_2 mpw5_submission_0/outd_0/InputSignal io_analog[3] io_analog[3] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12322 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12323 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12324 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12325 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12326 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12327 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12328 vccd1 mpw5_submission_1/isource_0/VM14D mpw5_submission_1/isource_0/VM12G mpw5_submission_1/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X12329 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12330 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12331 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12332 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12333 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12334 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12335 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12336 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X12337 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12338 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12339 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12340 a_429020_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12341 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12342 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12343 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12344 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12345 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12346 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12347 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12348 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12349 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12350 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12351 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12352 io_analog[5] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X12353 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12354 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12355 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12356 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12357 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12358 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12359 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12360 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12361 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12362 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12363 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12364 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12365 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D98 vssd1 io_analog[2] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X12366 a_442498_643680# mpw5_submission_0/cmirror_channel_0/I_in_channel vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12367 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12368 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12369 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12370 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12371 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12372 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12373 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12374 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_194220_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12375 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12376 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12377 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12378 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12379 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12380 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12381 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12382 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12383 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12384 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12385 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12386 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12387 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12388 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12389 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12390 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12391 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12392 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12393 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12394 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12395 mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X12396 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12397 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12398 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12399 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12400 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12401 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12402 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12403 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12404 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12405 a_427670_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12406 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12407 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12408 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X12409 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12410 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12411 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12412 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12413 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12414 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12415 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12416 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12417 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12418 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12419 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12420 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12421 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12422 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12423 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12424 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12425 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12426 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12427 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12428 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12429 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12430 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12431 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12432 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12433 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12434 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X12435 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12436 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12437 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12438 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12439 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12440 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12441 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12442 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12443 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12444 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12445 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12446 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12447 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12448 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12449 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12450 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X12451 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12452 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12453 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12454 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12455 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12456 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12457 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12458 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12459 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12460 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12461 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12462 a_184770_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12463 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12464 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12465 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12466 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12467 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12468 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12469 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12470 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12471 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12472 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12473 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12474 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12475 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12476 vssd1 vccd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X12477 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12478 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12479 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12480 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12481 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12482 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12483 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12484 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12485 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12486 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12487 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12488 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12489 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12490 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12491 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12492 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12493 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12494 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12495 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12496 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12497 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12498 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12499 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12500 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12501 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12502 vssd1 mpw5_submission_1/isource_0/VM11D a_181958_664870# vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X12503 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12504 a_430370_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12505 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12506 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12507 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12508 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12509 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12510 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12511 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12512 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12513 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12514 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12515 vccd1 io_analog[0] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X12516 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12517 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12518 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12519 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12520 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12521 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12522 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12523 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12524 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12525 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12526 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12527 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12528 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12529 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12530 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12531 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12532 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12533 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12534 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12535 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12536 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12537 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12538 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12539 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12540 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12541 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12542 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12543 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X12544 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12545 a_189936_658659# mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM8D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X12546 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12547 vssd1 mpw5_submission_0/cmirror_channel_0/I_in_channel a_441658_643680# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12548 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12549 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12550 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12551 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12552 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12553 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12554 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12555 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12556 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12557 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12558 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12559 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_184770_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12560 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12561 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12562 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_195570_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12563 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12564 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12565 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12566 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12567 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12568 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12569 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12570 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12571 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X12572 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12573 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12574 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12575 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12576 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12577 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12578 mpw5_submission_0/outd_0/InputSignal io_analog[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12579 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_190170_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12580 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12581 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12582 mpw5_submission_1/outd_0/V_da2_P vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X12583 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12584 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12585 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12586 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12587 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12588 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12589 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12590 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12591 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12592 a_441920_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12593 mpw5_submission_1/outd_0/InputSignal io_analog[6] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12594 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12595 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12596 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12597 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12598 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12599 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12600 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12601 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12602 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12603 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12604 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12605 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12606 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12607 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12608 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12609 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12610 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12611 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12612 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12613 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12614 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12615 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12616 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12617 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12618 a_200618_647480# mpw5_submission_1/cmirror_channel_0/I_in_channel vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12619 a_430136_648079# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X12620 mpw5_submission_1/outd_0/InputSignal io_analog[6] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12621 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12622 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12623 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12624 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12625 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12626 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12627 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12628 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12629 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12630 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12631 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_191520_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12632 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12633 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12634 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12635 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12636 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12637 a_435770_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12638 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12639 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12640 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12641 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12642 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12643 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12644 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12645 a_188820_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12646 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12647 mpw5_submission_0/isource_0/VM3D a_411216_644902# mpw5_submission_0/isource_0/VM22D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X12648 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12649 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12650 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12651 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12652 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12653 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12654 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12655 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12656 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12657 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12658 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12659 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12660 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12661 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12662 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12663 vssd1 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM5D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12664 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12665 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12666 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12667 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12668 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12669 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12670 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12671 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12672 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12673 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12674 vssd1 mpw5_submission_0/cmirror_channel_0/I_in_channel a_442498_643680# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12675 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12676 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12677 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12678 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12679 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12680 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12681 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12682 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12683 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12684 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12685 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12686 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12687 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12688 mpw5_submission_1/tia_core_0/VM36D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM39D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12689 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12690 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12691 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12692 mpw5_submission_1/tia_core_0/VM36D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM39D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12693 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12694 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12695 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12696 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12697 a_187470_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12698 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12699 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12700 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12701 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12702 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12703 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12704 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12705 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12706 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12707 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12708 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12709 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12710 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12711 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12712 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12713 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12714 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12715 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12716 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12717 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12718 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12719 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12720 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_464438_656600# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12721 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12722 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12723 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12724 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12725 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12726 a_440818_643680# mpw5_submission_0/cmirror_channel_0/I_in_channel vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12727 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12728 a_201458_647480# mpw5_submission_1/cmirror_channel_0/I_in_channel a_201520_649146# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12729 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12730 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12731 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12732 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12733 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12734 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12735 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12736 a_187976_652606# a_188506_655038# vssd1 sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X12737 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12738 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12739 a_433070_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12740 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12741 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12742 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12743 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12744 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12745 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12746 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12747 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12748 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12749 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12750 a_186120_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12751 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12752 mpw5_submission_1/outd_0/InputSignal io_analog[6] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12753 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12754 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12755 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12756 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12757 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12758 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12759 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12760 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12761 io_analog[2] mpw5_submission_0/eigth_mirror_0/I_In a_433070_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12762 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12763 io_analog[3] mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM5D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12764 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12765 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12766 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12767 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12768 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12769 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12770 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12771 vssd1 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM5D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12772 mpw5_submission_1/outd_0/InputSignal io_analog[6] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12773 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12774 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12775 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12776 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12777 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12778 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12779 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12780 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12781 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12782 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12783 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12784 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12785 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_658659# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X12786 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12787 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12788 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12789 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12790 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12791 a_181958_664870# mpw5_submission_1/isource_0/VM11D vssd1 vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X12792 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12793 a_189936_651879# mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM14D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X12794 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12795 vccd1 mpw5_submission_0/tia_core_0/VM40D sky130_fd_pr__cap_mim_m3_2 l=1.8e+07u w=2.5e+07u
X12796 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12797 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12798 a_189936_658659# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X12799 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12800 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12801 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12802 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12803 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12804 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12805 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12806 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12807 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12808 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12809 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12810 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12811 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12812 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12813 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X12814 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12815 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12816 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12817 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12818 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12819 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12820 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12821 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12822 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12823 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12824 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12825 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12826 a_443570_645443# a_441720_645346# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12827 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12828 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12829 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12830 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12831 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12832 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12833 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12834 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12835 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12836 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12837 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12838 vccd1 io_analog[5] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X12839 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12840 a_441720_645346# mpw5_submission_0/cmirror_channel_0/I_in_channel a_441658_643680# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12841 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12842 vssd1 mpw5_submission_0/isource_0/VM11D a_422158_661070# vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X12843 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12844 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12845 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12846 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12847 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12848 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12849 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12850 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12851 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12852 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D99 vssd1 io_analog[8] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X12853 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12854 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12855 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12856 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12857 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12858 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12859 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12860 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12861 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12862 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12863 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12864 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12865 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12866 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12867 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12868 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12869 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12870 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12871 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12872 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12873 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12874 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12875 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12876 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12877 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_654859# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X12878 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12879 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12880 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12881 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12882 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12883 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12884 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12885 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12886 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12887 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12888 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12889 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12890 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X12891 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12892 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12893 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12894 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12895 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12896 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12897 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D100 vssd1 io_analog[7] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X12898 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12899 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12900 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12901 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12902 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12903 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12904 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12905 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12906 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12907 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12908 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12909 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12910 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12911 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12912 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12913 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12914 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12915 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12916 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12917 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12918 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12919 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12920 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12921 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12922 mpw5_submission_0/tia_core_0/Out_2 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12923 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12924 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12925 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12926 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X12927 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12928 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12929 mpw5_submission_0/outd_0/InputSignal io_analog[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12930 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12931 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12932 mpw5_submission_1/tia_core_0/VM5D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 io_analog[6] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12933 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12934 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12935 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12936 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12937 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12938 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12939 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12940 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12941 a_427670_636823# mpw5_submission_0/eigth_mirror_0/I_In mpw5_submission_0/eigth_mirror_0/I_out_5 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12942 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12943 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12944 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12945 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12946 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12947 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12948 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12949 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12950 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12951 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12952 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12953 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12954 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12955 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12956 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12957 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12958 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12959 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12960 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12961 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12962 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12963 vccd1 io_analog[5] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X12964 mpw5_submission_1/tia_core_0/Out_2 mpw5_submission_1/outd_0/InputSignal io_analog[6] io_analog[6] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12965 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12966 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12967 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12968 a_443850_641883# a_441720_645346# mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12969 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12970 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12971 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12972 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12973 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12974 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12975 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12976 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12977 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12978 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12979 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12980 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12981 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12982 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12983 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12984 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12985 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12986 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12987 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12988 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12989 a_426320_636823# mpw5_submission_0/eigth_mirror_0/I_In mpw5_submission_0/eigth_mirror_0/I_out_6 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12990 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12991 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12992 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12993 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12994 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12995 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12996 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12997 a_203650_645683# a_201520_649146# mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12998 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12999 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13000 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13001 mpw5_submission_0/outd_0/InputSignal io_analog[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13002 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13003 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13004 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13005 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13006 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13007 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13008 vccd1 io_analog[5] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X13009 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13010 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13011 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13012 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13013 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13014 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13015 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13016 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13017 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13018 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13019 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13020 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13021 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13022 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13023 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13024 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13025 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13026 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X13027 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13028 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13029 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13030 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13031 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13032 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13033 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13034 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13035 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13036 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM6D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13037 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13038 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13039 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13040 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13041 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13042 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D101 io_analog[1] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X13043 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D102 io_analog[0] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X13044 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13045 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13046 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13047 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13048 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13049 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13050 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13051 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13052 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13053 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13054 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13055 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13056 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13057 a_411216_644902# mpw5_submission_0/isource_0/VM22D mpw5_submission_0/eigth_mirror_0/I_In vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X13058 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13059 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13060 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13061 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13062 io_analog[1] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X13063 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13064 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13065 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13066 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13067 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13068 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13069 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X13070 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13071 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13072 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13073 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13074 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13075 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13076 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13077 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13078 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13079 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13080 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13081 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13082 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13083 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13084 a_430136_648079# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X13085 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13086 vccd1 io_analog[3] mpw5_submission_0/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13087 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13088 io_analog[3] mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/tia_core_0/Out_2 io_analog[3] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13089 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13090 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13091 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13092 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13093 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13094 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13095 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13096 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13097 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13098 a_427670_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13099 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13100 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13101 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13102 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13103 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13104 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13105 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13106 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13107 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13108 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13109 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13110 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13111 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13112 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13113 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13114 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13115 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13116 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13117 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13118 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13119 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13120 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13121 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13122 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13123 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13124 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13125 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13126 mpw5_submission_0/tia_core_0/VM31D vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13127 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13128 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13129 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13130 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13131 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13132 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13133 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13134 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13135 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13136 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13137 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13138 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13139 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13140 vccd1 mpw5_submission_0/isource_0/VM14D mpw5_submission_0/isource_0/VM12G mpw5_submission_0/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X13141 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13142 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X13143 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13144 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13145 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13146 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13147 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13148 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13149 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13150 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13151 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13152 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13153 a_422158_661070# mpw5_submission_0/isource_0/VM11D vssd1 vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X13154 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13155 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13156 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X13157 a_426320_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13158 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13159 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13160 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13161 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13162 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13163 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13164 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13165 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13166 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13167 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13168 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D103 vssd1 io_analog[1] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X13169 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13170 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13171 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13172 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13173 a_430136_648079# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X13174 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13175 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13176 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13177 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13178 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13179 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13180 mpw5_submission_0/tia_core_0/Out_2 mpw5_submission_0/outd_0/InputSignal io_analog[3] io_analog[3] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13181 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13182 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13183 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13184 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13185 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13186 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13187 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13188 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13189 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
D104 io_analog[2] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X13190 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13191 io_analog[1] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X13192 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13193 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13194 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13195 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13196 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13197 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13198 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13199 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13200 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13201 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13202 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13203 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13204 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13205 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13206 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13207 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13208 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13209 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13210 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13211 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13212 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13213 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/InputRef mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13214 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13215 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13216 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13217 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13218 a_424970_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13219 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13220 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13221 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13222 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13223 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13224 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13225 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13226 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13227 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13228 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13229 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_433070_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13230 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13231 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13232 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13233 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13234 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_430370_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13235 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13236 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13237 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13238 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13239 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13240 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13241 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13242 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13243 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13244 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13245 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13246 vssd1 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM6D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13247 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13248 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_433070_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13249 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13250 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13251 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13252 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13253 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13254 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X13255 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13256 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13257 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13258 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13259 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13260 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13261 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13262 a_203650_645683# a_201520_649146# mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13263 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13264 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13265 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13266 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13267 vccd1 io_analog[4] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X13268 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13269 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13270 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13271 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X13272 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13273 vccd1 mpw5_submission_0/isource_0/VM8D sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X13274 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13275 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13276 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13277 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM2D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X13278 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13279 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13280 io_analog[1] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X13281 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13282 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13283 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13284 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13285 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13286 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13287 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13288 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13289 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13290 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_431720_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13291 a_443850_641883# a_441720_645346# mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13292 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13293 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13294 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13295 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13296 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13297 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13298 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13299 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
R5 vssd1 io_clamp_low[1] sky130_fd_pr__res_generic_m3 w=1.1e+07u l=250000u
X13300 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_434420_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13301 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13302 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13303 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13304 vccd1 io_analog[4] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X13305 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13306 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13307 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13308 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13309 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13310 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_187470_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13311 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13312 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13313 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13314 vssd1 io_analog[7] mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=1e+06u
X13315 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13316 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13317 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13318 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13319 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13320 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13321 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13322 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13323 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13324 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13325 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13326 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13327 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13328 vccd1 mpw5_submission_1/isource_0/VM11D a_181958_664870# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X13329 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13330 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13331 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13332 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13333 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13334 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13335 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13336 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13337 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13338 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13339 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13340 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13341 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13342 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13343 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13344 io_analog[4] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X13345 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13346 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13347 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13348 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13349 mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X13350 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13351 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X13352 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D105 vssd1 io_analog[3] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X13353 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13354 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13355 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13356 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13357 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13358 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13359 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13360 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13361 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13362 vssd1 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM6D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13363 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13364 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13365 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13366 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13367 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM31D mpw5_submission_0/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13368 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13369 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13370 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13371 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13372 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13373 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13374 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13375 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13376 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13377 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13378 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D106 io_analog[8] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X13379 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13380 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X13381 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13382 vssd1 a_188506_655038# vssd1 sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X13383 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X13384 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X13385 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13386 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13387 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13388 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13389 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13390 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13391 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13392 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13393 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13394 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13395 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13396 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13397 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13398 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13399 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13400 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13401 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13402 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13403 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13404 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13405 mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/InputRef mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13406 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13407 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13408 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13409 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13410 io_analog[3] mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/tia_core_0/Out_2 io_analog[3] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13411 mpw5_submission_0/isource_0/VM3D a_411216_644902# mpw5_submission_0/isource_0/VM22D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X13412 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13413 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13414 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13415 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13416 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13417 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13418 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13419 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13420 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13421 a_429020_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13422 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13423 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13424 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13425 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13426 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13427 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13428 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13429 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13430 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13431 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13432 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13433 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13434 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13435 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13436 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13437 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13438 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13439 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13440 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13441 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13442 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13443 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13444 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13445 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13446 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13447 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13448 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13449 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13450 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13451 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13452 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13453 vssd1 io_analog[7] mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13454 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13455 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM36D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13456 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13457 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13458 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13459 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13460 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13461 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13462 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13463 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13464 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13465 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13466 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13467 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13468 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13469 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13470 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13471 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13472 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13473 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13474 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13475 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13476 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13477 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13478 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13479 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13480 a_192870_640623# mpw5_submission_1/eigth_mirror_0/I_In mpw5_submission_1/eigth_mirror_0/I_out_1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13481 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13482 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13483 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13484 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13485 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13486 a_427670_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13487 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13488 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13489 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13490 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13491 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13492 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13493 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13494 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_464438_656600# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13495 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X13496 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X13497 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13498 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13499 mpw5_submission_1/isource_0/VM3G a_184186_655038# vssd1 sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X13500 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13501 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13502 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13503 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13504 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13505 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13506 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13507 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13508 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13509 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13510 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13511 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13512 a_424970_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13513 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13514 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13515 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13516 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13517 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13518 a_443570_645443# a_441720_645346# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13519 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13520 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13521 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13522 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13523 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13524 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13525 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13526 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13527 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13528 mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__cap_var_lvt pd=0u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X13529 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13530 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13531 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13532 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13533 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13534 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13535 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13536 a_191520_640623# mpw5_submission_1/eigth_mirror_0/I_In mpw5_submission_1/eigth_mirror_0/I_out_2 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13537 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13538 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13539 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13540 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13541 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13542 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13543 a_201720_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13544 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13545 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13546 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13547 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_190170_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13548 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13549 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13550 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D107 vssd1 io_analog[2] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X13551 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13552 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13553 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13554 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13555 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13556 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13557 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13558 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13559 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13560 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13561 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13562 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13563 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13564 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13565 a_441920_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13566 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13567 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13568 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13569 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13570 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13571 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13572 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13573 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13574 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13575 mpw5_submission_0/isource_0/VM3D a_411216_644902# mpw5_submission_0/isource_0/VM22D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X13576 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13577 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM31D mpw5_submission_0/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13578 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13579 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13580 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13581 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13582 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13583 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13584 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13585 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13586 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13587 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13588 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13589 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13590 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13591 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13592 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13593 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13594 vssd1 mpw5_submission_1/isource_0/VM11D a_181958_664870# vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X13595 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13596 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13597 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13598 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13599 mpw5_submission_1/tia_core_0/VM36D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13600 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13601 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13602 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13603 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13604 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13605 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13606 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D108 io_analog[1] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X13607 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_191520_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13608 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13609 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13610 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13611 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13612 vccd1 a_201520_649146# a_201720_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13613 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13614 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13615 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13616 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13617 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13618 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13619 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13620 vssd1 vccd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X13621 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13622 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13623 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13624 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13625 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13626 mpw5_submission_1/outd_0/InputSignal io_analog[6] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13627 vssd1 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM5D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13628 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13629 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13630 a_203370_649243# a_201520_649146# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13631 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13632 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13633 mpw5_submission_1/isource_0/VM3D a_171016_648702# mpw5_submission_1/isource_0/VM22D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X13634 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13635 mpw5_submission_0/isource_0/VM22D a_411216_644902# mpw5_submission_0/isource_0/VM3D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X13636 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13637 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13638 mpw5_submission_0/isource_0/VM22D a_411216_644902# mpw5_submission_0/isource_0/VM3D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X13639 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13640 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13641 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13642 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13643 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13644 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13645 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13646 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13647 mpw5_submission_1/tia_core_0/VM6D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13648 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13649 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13650 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13651 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13652 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13653 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13654 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13655 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_190170_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13656 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13657 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13658 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13659 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13660 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13661 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X13662 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13663 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13664 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13665 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13666 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13667 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13668 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13669 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13670 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13671 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13672 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13673 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13674 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13675 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13676 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13677 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13678 a_430136_648079# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X13679 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13680 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13681 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13682 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13683 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13684 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13685 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224238_660400# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13686 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13687 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13688 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13689 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13690 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13691 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13692 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13693 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13694 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13695 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13696 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X13697 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13698 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13699 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13700 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13701 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13702 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13703 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13704 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13705 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13706 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13707 mpw5_submission_1/outd_0/InputSignal io_analog[6] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13708 vccd1 mpw5_submission_1/tia_core_0/VM40D sky130_fd_pr__cap_mim_m3_2 l=1.8e+07u w=2.5e+07u
X13709 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13710 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13711 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13712 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13713 a_191520_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13714 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13715 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13716 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13717 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13718 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13719 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13720 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13721 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13722 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13723 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13724 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13725 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13726 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13727 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13728 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13729 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13730 mpw5_submission_1/outd_0/InputSignal io_analog[6] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13731 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13732 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13733 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13734 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13735 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13736 io_analog[6] mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM5D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13737 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13738 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13739 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13740 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13741 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D109 vssd1 io_analog[8] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X13742 vssd1 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM5D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13743 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13744 mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X13745 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13746 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13747 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13748 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13749 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13750 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13751 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13752 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13753 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13754 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13755 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13756 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13757 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13758 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13759 io_analog[0] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X13760 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13761 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13762 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13763 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13764 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13765 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13766 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13767 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13768 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13769 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13770 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13771 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13772 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13773 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_660919# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X13774 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13775 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13776 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13777 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13778 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13779 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13780 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM31D mpw5_submission_1/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13781 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13782 a_191520_640623# mpw5_submission_1/eigth_mirror_0/I_In mpw5_submission_1/eigth_mirror_0/I_out_2 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13783 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13784 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13785 vccd1 mpw5_submission_0/outd_0/V_da2_N vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X13786 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13787 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13788 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13789 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X13790 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13791 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13792 mpw5_submission_0/isource_0/VM22D a_411216_644902# mpw5_submission_0/isource_0/VM3D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X13793 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13794 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13795 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13796 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13797 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13798 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13799 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13800 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13801 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13802 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13803 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_658659# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X13804 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13805 vccd1 io_analog[0] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X13806 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13807 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13808 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13809 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13810 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13811 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13812 a_187976_652606# a_187446_655038# vssd1 sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X13813 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13814 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13815 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13816 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13817 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13818 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13819 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13820 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13821 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13822 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13823 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13824 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13825 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13826 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X13827 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13828 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13829 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13830 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13831 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13832 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13833 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13834 mpw5_submission_0/tia_core_0/VM5D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 io_analog[3] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13835 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13836 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13837 vccd1 vssd1 mpw5_submission_0/tia_core_0/VM31D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13838 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13839 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13840 mpw5_submission_1/outd_0/V_da2_N vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X13841 mpw5_submission_1/tia_core_0/VM6D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13842 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X13843 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13844 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13845 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13846 vccd1 io_analog[5] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X13847 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13848 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13849 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13850 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13851 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X13852 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13853 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13854 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X13855 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13856 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13857 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13858 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13859 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13860 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13861 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13862 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13863 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13864 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13865 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13866 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13867 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13868 mpw5_submission_0/eigth_mirror_0/I_In mpw5_submission_0/isource_0/VM22D a_411216_644902# vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X13869 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13870 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13871 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13872 mpw5_submission_1/tia_core_0/Out_2 mpw5_submission_1/outd_0/InputSignal io_analog[6] io_analog[6] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13873 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13874 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13875 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13876 io_analog[2] mpw5_submission_0/eigth_mirror_0/I_In a_433070_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13877 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13878 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13879 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13880 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13881 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13882 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13883 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13884 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13885 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13886 io_analog[6] mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/tia_core_0/Out_2 io_analog[6] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13887 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13888 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13889 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13890 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13891 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13892 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13893 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13894 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13895 mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X13896 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13897 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13898 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13899 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13900 mpw5_submission_0/tia_core_0/VM31D mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13901 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13902 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13903 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13904 mpw5_submission_0/outd_0/InputSignal io_analog[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13905 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13906 mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__cap_var_lvt pd=0u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X13907 mpw5_submission_1/tia_core_0/Out_2 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13908 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13909 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13910 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13911 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13912 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13913 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13914 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D110 io_analog[7] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X13915 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13916 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13917 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13918 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13919 a_181958_664870# mpw5_submission_1/isource_0/VM11D vssd1 vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X13920 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13921 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13922 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13923 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13924 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13925 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13926 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13927 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13928 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13929 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13930 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13931 mpw5_submission_0/isource_0/VM12G mpw5_submission_0/isource_0/VM14D vccd1 mpw5_submission_0/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X13932 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13933 mpw5_submission_0/isource_0/VM12G mpw5_submission_0/isource_0/VM14D vccd1 mpw5_submission_0/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X13934 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13935 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13936 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13937 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13938 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13939 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13940 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13941 a_443570_645443# a_441720_645346# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13942 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13943 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13944 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13945 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13946 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13947 vssd1 vccd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X13948 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13949 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13950 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13951 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13952 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13953 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X13954 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13955 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13956 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13957 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13958 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13959 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13960 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13961 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13962 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13963 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13964 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13965 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X13966 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13967 vssd1 mpw5_submission_0/isource_0/VM11D a_422158_661070# vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X13968 a_194220_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13969 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13970 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13971 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13972 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13973 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13974 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13975 a_430136_657119# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X13976 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13977 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13978 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13979 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13980 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13981 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13982 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13983 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13984 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13985 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13986 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13987 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D111 io_analog[3] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X13988 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13989 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13990 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13991 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13992 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13993 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_427670_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13994 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13995 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X13996 vccd1 io_analog[4] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X13997 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13998 mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/InputRef mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13999 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14000 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14001 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14002 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14003 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14004 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14005 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14006 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14007 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14008 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14009 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14010 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14011 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14012 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14013 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14014 mpw5_submission_0/tia_core_0/VM36D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14015 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14016 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14017 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14018 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14019 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14020 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14021 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14022 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14023 a_203650_645683# a_201520_649146# mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14024 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14025 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14026 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14027 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14028 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14029 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14030 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14031 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14032 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14033 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14034 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14035 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14036 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14037 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14038 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14039 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14040 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14041 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14042 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14043 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14044 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14045 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14046 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14047 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14048 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14049 a_200618_647480# mpw5_submission_1/cmirror_channel_0/I_in_channel vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14050 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14051 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14052 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14053 io_analog[1] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X14054 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14055 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14056 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14057 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X14058 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14059 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14060 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14061 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14062 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14063 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14064 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14065 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14066 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14067 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14068 vssd1 vccd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X14069 vccd1 mpw5_submission_1/outd_0/V_da2_P vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X14070 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14071 mpw5_submission_0/outd_0/InputSignal io_analog[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14072 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14073 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14074 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14075 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14076 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X14077 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14078 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14079 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X14080 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14081 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14082 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14083 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14084 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14085 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14086 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14087 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14088 io_analog[6] mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/tia_core_0/Out_2 io_analog[6] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14089 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14090 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14091 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14092 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14093 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14094 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14095 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14096 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14097 a_411216_644902# mpw5_submission_0/isource_0/VM22D mpw5_submission_0/eigth_mirror_0/I_In vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X14098 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14099 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14100 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14101 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14102 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14103 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14104 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14105 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14106 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14107 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14108 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14109 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14110 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14111 mpw5_submission_1/tia_core_0/Out_2 mpw5_submission_1/outd_0/InputSignal io_analog[6] io_analog[6] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14112 a_201720_649243# a_201520_649146# a_201520_649146# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14113 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14114 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14115 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14116 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14117 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14118 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14119 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14120 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14121 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14122 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14123 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14124 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14125 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14126 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14127 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14128 a_441658_643680# mpw5_submission_0/cmirror_channel_0/I_in_channel vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14129 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14130 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14131 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14132 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14133 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14134 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14135 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14136 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14137 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14138 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14139 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14140 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14141 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14142 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14143 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14144 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14145 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14146 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14147 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14148 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14149 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14150 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14151 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14152 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14153 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14154 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14155 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14156 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14157 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14158 mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/InputRef mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14159 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14160 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14161 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14162 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14163 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14164 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14165 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14166 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14167 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14168 mpw5_submission_0/eigth_mirror_0/I_In mpw5_submission_0/isource_0/VM22D a_411216_644902# vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X14169 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14170 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_184770_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14171 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14172 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14173 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14174 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_195570_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14175 vccd1 mpw5_submission_0/tia_core_0/VM28D sky130_fd_pr__cap_mim_m3_2 l=1.8e+07u w=2.5e+07u
X14176 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14177 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14178 vccd1 mpw5_submission_0/isource_0/VM14D mpw5_submission_0/isource_0/VM12G mpw5_submission_0/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X14179 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14180 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14181 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14182 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM2D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X14183 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14184 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14185 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14186 a_430136_648079# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X14187 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14188 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14189 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14190 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14191 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14192 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14193 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14194 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/InputRef mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14195 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14196 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14197 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/InputRef mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14198 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14199 io_analog[6] mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/tia_core_0/Out_2 io_analog[6] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14200 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14201 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14202 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14203 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14204 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14205 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X14206 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14207 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14208 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14209 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14210 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14211 mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__cap_var_lvt pd=0u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X14212 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14213 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14214 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14215 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14216 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14217 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14218 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14219 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14220 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14221 mpw5_submission_0/tia_core_0/Out_2 mpw5_submission_0/outd_0/InputSignal io_analog[3] io_analog[3] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14222 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14223 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_186120_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14224 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14225 vccd1 vssd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X14226 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14227 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14228 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14229 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14230 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14231 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14232 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14233 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14234 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_194220_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14235 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14236 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14237 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14238 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14239 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14240 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14241 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14242 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14243 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14244 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14245 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14246 a_187470_640623# mpw5_submission_1/eigth_mirror_0/I_In mpw5_submission_1/eigth_mirror_0/I_out_5 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14247 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14248 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14249 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 io_analog[7] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14250 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14251 mpw5_submission_1/tia_core_0/VM36D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM39D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14252 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_433070_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14253 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14254 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14255 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14256 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14257 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14258 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14259 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14260 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_191520_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14261 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14262 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14263 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14264 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14265 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14266 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14267 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14268 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14269 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14270 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14271 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14272 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14273 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14274 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14275 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14276 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14277 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14278 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14279 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14280 a_430136_648079# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X14281 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14282 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14283 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14284 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14285 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14286 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14287 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14288 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14289 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14290 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14291 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14292 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14293 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14294 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
R6 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA sky130_fd_pr__res_generic_m3 w=1.5e+06u l=500000u
X14295 mpw5_submission_1/eigth_mirror_0/I_out_1 mpw5_submission_1/eigth_mirror_0/I_In a_192870_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14296 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14297 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14298 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14299 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14300 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14301 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14302 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14303 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14304 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14305 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14306 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14307 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14308 mpw5_submission_0/outd_0/V_da2_P vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X14309 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14310 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14311 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14312 a_411216_644902# mpw5_submission_0/isource_0/VM22D mpw5_submission_0/eigth_mirror_0/I_In vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X14313 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14314 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_434420_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14315 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14316 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D112 io_analog[7] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X14317 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14318 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14319 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14320 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_187470_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14321 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14322 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14323 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14324 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14325 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14326 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14327 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14328 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14329 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14330 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14331 mpw5_submission_0/tia_core_0/Out_2 mpw5_submission_0/outd_0/InputSignal io_analog[3] io_analog[3] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14332 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14333 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14334 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14335 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X14336 io_analog[1] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X14337 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14338 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14339 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14340 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14341 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14342 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14343 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14344 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14345 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14346 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14347 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14348 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14349 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14350 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14351 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_433070_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14352 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14353 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14354 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14355 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_430370_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14356 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14357 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14358 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14359 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14360 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14361 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14362 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14363 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14364 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14365 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14366 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14367 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14368 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14369 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14370 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14371 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14372 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14373 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14374 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14375 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14376 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14377 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14378 vccd1 io_analog[1] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X14379 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14380 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14381 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14382 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14383 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14384 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14385 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14386 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14387 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14388 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14389 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14390 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14391 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14392 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14393 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14394 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14395 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14396 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14397 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14398 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14399 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14400 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14401 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14402 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14403 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14404 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14405 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14406 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14407 a_171016_648702# mpw5_submission_1/isource_0/VM22D mpw5_submission_1/eigth_mirror_0/I_In vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X14408 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14409 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14410 a_429020_636823# mpw5_submission_0/eigth_mirror_0/I_In mpw5_submission_0/eigth_mirror_0/I_out_4 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14411 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14412 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_431720_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14413 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14414 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14415 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14416 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14417 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14418 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14419 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_184770_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14420 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14421 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14422 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14423 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14424 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14425 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X14426 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14427 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14428 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14429 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14430 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14431 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14432 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14433 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14434 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14435 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14436 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14437 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14438 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14439 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14440 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14441 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14442 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14443 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14444 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14445 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14446 mpw5_submission_0/cmirror_channel_0/I_in_channel mpw5_submission_0/eigth_mirror_0/I_In a_434420_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14447 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14448 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14449 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14450 io_analog[0] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X14451 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14452 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14453 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14454 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14455 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14456 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14457 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14458 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14459 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14460 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14461 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14462 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14463 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14464 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14465 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14466 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14467 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14468 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14469 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14470 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14471 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14472 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14473 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14474 vccd1 mpw5_submission_1/tia_core_0/VM28D sky130_fd_pr__cap_mim_m3_2 l=1.8e+07u w=2.5e+07u
X14475 a_186120_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14476 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14477 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14478 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14479 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14480 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14481 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14482 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14483 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14484 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14485 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14486 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14487 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14488 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14489 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14490 a_187470_640623# mpw5_submission_1/eigth_mirror_0/I_In mpw5_submission_1/eigth_mirror_0/I_out_5 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14491 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14492 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14493 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14494 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14495 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14496 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14497 a_194220_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14498 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14499 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14500 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14501 a_424970_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14502 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14503 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14504 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14505 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14506 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14507 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14508 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14509 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14510 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14511 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14512 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14513 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14514 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14515 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14516 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14517 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14518 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14519 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X14520 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14521 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14522 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14523 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14524 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14525 vccd1 vssd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X14526 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14527 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14528 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14529 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14530 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14531 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14532 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14533 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14534 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14535 mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X14536 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14537 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14538 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14539 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14540 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14541 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14542 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14543 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14544 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14545 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14546 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14547 a_186120_640623# mpw5_submission_1/eigth_mirror_0/I_In mpw5_submission_1/eigth_mirror_0/I_out_6 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14548 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14549 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14550 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14551 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14552 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14553 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14554 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14555 io_analog[3] mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/tia_core_0/Out_2 io_analog[3] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14556 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14557 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14558 a_192870_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14559 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14560 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14561 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14562 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14563 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14564 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14565 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14566 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14567 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14568 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14569 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14570 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14571 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14572 mpw5_submission_1/tia_core_0/VM6D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14573 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14574 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14575 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14576 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14577 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14578 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14579 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14580 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14581 a_442498_643680# mpw5_submission_0/cmirror_channel_0/I_in_channel vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14582 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14583 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14584 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14585 mpw5_submission_1/tia_core_0/VM31D mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14586 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14587 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14588 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14589 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14590 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14591 vssd1 vccd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X14592 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14593 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14594 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14595 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14596 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14597 vccd1 a_441720_645346# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X14598 mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__cap_var_lvt pd=0u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X14599 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14600 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14601 a_430136_645809# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X14602 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14603 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14604 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14605 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14606 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14607 vccd1 io_analog[1] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X14608 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14609 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14610 a_430136_648079# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X14611 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14612 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14613 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14614 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14615 io_analog[3] mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_0/tia_core_0/VM5D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14616 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM6D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14617 io_analog[5] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X14618 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14619 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14620 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14621 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14622 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14623 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14624 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14625 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14626 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14627 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14628 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14629 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14630 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14631 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14632 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14633 mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM9D mpw5_submission_0/isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X14634 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14635 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14636 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14637 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14638 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14639 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14640 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14641 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14642 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14643 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14644 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14645 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14646 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14647 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D113 vssd1 io_analog[3] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X14648 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14649 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14650 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14651 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14652 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14653 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14654 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14655 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14656 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14657 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14658 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14659 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14660 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14661 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14662 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14663 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14664 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14665 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14666 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14667 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14668 vccd1 mpw5_submission_1/isource_0/VM14D mpw5_submission_1/isource_0/VM12G mpw5_submission_1/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X14669 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14670 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D114 vssd1 io_analog[1] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X14671 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14672 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14673 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14674 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14675 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14676 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X14677 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14678 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14679 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X14680 vccd1 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14681 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14682 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14683 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14684 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14685 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM31D mpw5_submission_0/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14686 mpw5_submission_1/tia_core_0/VM31D vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14687 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14688 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14689 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14690 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14691 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14692 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14693 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14694 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14695 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14696 a_203650_645683# a_201520_649146# mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14697 a_189936_651879# mpw5_submission_1/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X14698 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14699 vccd1 mpw5_submission_0/isource_0/VM14D mpw5_submission_0/isource_0/VM12G mpw5_submission_0/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X14700 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14701 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14702 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14703 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14704 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14705 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14706 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14707 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14708 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14709 vssd1 mpw5_submission_1/isource_0/VM11D a_181958_664870# vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X14710 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14711 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14712 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14713 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14714 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14715 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14716 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14717 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14718 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14719 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14720 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14721 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14722 a_189936_660919# mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM9D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X14723 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14724 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14725 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14726 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14727 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14728 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14729 vssd1 mpw5_submission_0/cmirror_channel_0/I_in_channel a_441658_643680# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14730 a_430136_648079# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X14731 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14732 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14733 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14734 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14735 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14736 mpw5_submission_1/outd_0/InputSignal io_analog[6] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14737 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14738 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D115 io_analog[1] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X14739 vccd1 mpw5_submission_1/isource_0/VM8D a_189936_651879# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X14740 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14741 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14742 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14743 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14744 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14745 vccd1 io_analog[0] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X14746 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14747 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14748 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14749 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14750 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14751 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14752 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14753 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14754 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14755 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14756 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14757 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14758 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14759 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14760 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14761 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14762 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14763 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14764 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14765 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14766 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14767 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14768 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/InputRef mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14769 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14770 mpw5_submission_0/tia_core_0/VM31D mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14771 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14772 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14773 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14774 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14775 vccd1 io_analog[1] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X14776 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14777 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14778 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14779 mpw5_submission_0/tia_core_0/VM31D vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14780 a_202298_647480# mpw5_submission_1/cmirror_channel_0/I_in_channel vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14781 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14782 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14783 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14784 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14785 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14786 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14787 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14788 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14789 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14790 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14791 mpw5_submission_1/tia_core_0/VM28D io_analog[6] mpw5_submission_1/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14792 mpw5_submission_1/tia_core_0/VM5D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 io_analog[6] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14793 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14794 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14795 a_195570_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14796 mpw5_submission_1/tia_core_0/VM5D mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 io_analog[6] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14797 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X14798 vssd1 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM6D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14799 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14800 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14801 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14802 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14803 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14804 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14805 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14806 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14807 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14808 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14809 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14810 mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14811 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14812 a_430136_648079# mpw5_submission_0/isource_0/VM8D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X14813 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14814 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14815 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14816 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14817 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14818 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14819 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14820 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14821 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14822 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14823 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14824 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14825 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X14826 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14827 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14828 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14829 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14830 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14831 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14832 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14833 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14834 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14835 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14836 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14837 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14838 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14839 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14840 vccd1 io_analog[0] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X14841 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14842 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14843 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14844 mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14845 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14846 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14847 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14848 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14849 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14850 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14851 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14852 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14853 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14854 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14855 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14856 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14857 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14858 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14859 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14860 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14861 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14862 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14863 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14864 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14865 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14866 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14867 vccd1 a_441720_645346# a_443570_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14868 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14869 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14870 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14871 mpw5_submission_1/outd_0/V_da2_N vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X14872 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=1e+06u
X14873 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14874 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14875 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14876 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14877 mpw5_submission_0/eigth_mirror_0/I_In mpw5_submission_0/isource_0/VM22D a_411216_644902# vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X14878 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14879 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14880 mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__cap_var_lvt pd=0u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X14881 a_430136_648079# mpw5_submission_0/isource_0/VM8D mpw5_submission_0/isource_0/VM14D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X14882 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14883 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14884 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14885 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14886 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14887 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14888 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14889 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14890 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14891 io_analog[4] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X14892 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14893 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14894 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14895 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14896 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14897 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14898 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14899 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14900 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14901 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14902 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14903 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14904 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X14905 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X14906 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14907 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14908 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14909 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14910 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14911 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14912 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14913 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14914 a_201520_649146# a_201520_649146# a_201720_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14915 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14916 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14917 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14918 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14919 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D116 io_analog[7] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X14920 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14921 mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14922 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14923 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14924 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14925 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14926 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14927 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14928 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14929 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14930 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_431720_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14931 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14932 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14933 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14934 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14935 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14936 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14937 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14938 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14939 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14940 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14941 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14942 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14943 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14944 mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/InputRef mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14945 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14946 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14947 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14948 a_189936_651879# mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM14D vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X14949 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14950 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14951 a_411216_644902# mpw5_submission_0/isource_0/VM22D mpw5_submission_0/eigth_mirror_0/I_In vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X14952 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14953 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14954 mpw5_submission_1/isource_0/VM3D a_171016_648702# mpw5_submission_1/isource_0/VM22D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X14955 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14956 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14957 mpw5_submission_0/isource_0/VM22D a_411216_644902# mpw5_submission_0/isource_0/VM3D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X14958 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14959 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14960 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_187470_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14961 mpw5_submission_0/isource_0/VM12G mpw5_submission_0/isource_0/VM14D vccd1 mpw5_submission_0/isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X14962 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14963 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14964 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14965 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14966 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14967 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14968 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14969 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14970 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14971 vssd1 mpw5_submission_1/cmirror_channel_0/I_in_channel a_201458_647480# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14972 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14973 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14974 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14975 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14976 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14977 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14978 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14979 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14980 mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/InputRef mpw5_submission_1/outd_0/outd_stage1_0/isource_out mpw5_submission_1/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14981 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14982 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14983 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14984 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14985 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14986 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14987 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14988 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14989 vssd1 vccd1 sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X14990 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14991 mpw5_submission_0/tia_core_0/VM6D mpw5_submission_0/cmirror_channel_0/TIA_I_Bias1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14992 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14993 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14994 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14995 mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X14996 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14997 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14998 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14999 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15000 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15001 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15002 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15003 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15004 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15005 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15006 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15007 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15008 mpw5_submission_1/tia_core_0/Out_2 mpw5_submission_1/outd_0/InputSignal io_analog[6] io_analog[6] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15009 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15010 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15011 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15012 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15013 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15014 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15015 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15016 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15017 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15018 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15019 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15020 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15021 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15022 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15023 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15024 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_186120_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15025 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15026 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15027 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15028 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15029 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15030 mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM31D mpw5_submission_0/tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15031 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15032 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15033 a_203370_649243# a_201520_649146# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15034 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15035 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15036 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15037 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15038 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15039 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15040 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15041 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15042 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15043 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15044 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15045 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15046 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15047 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15048 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15049 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15050 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15051 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15052 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15053 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15054 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15055 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15056 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15057 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15058 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15059 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15060 mpw5_submission_0/outd_0/InputSignal io_analog[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15061 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15062 vssd1 mpw5_submission_0/isource_0/VM12G mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X15063 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15064 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15065 mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15066 a_441920_645443# a_441720_645346# a_441720_645346# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15067 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15068 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15069 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15070 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15071 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15072 mpw5_submission_0/outd_0/InputRef mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15073 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15074 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15075 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15076 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15077 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15078 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15079 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15080 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15081 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15082 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15083 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15084 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15085 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15086 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15087 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15088 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15089 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X15090 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15091 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15092 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15093 a_203370_649243# a_201520_649146# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15094 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15095 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15096 vccd1 io_analog[0] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X15097 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15098 vccd1 io_analog[6] mpw5_submission_1/outd_0/InputSignal vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15099 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15100 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15101 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15102 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15103 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15104 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15105 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15106 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15107 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15108 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15109 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15110 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15111 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15112 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15113 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15114 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15115 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15116 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15117 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_427670_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15118 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15119 mpw5_submission_0/isource_0/VM22D a_411216_644902# mpw5_submission_0/isource_0/VM3D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X15120 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15121 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15122 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15123 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15124 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15125 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15126 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15127 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15128 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15129 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15130 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15131 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15132 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15133 io_analog[3] mpw5_submission_0/outd_0/InputSignal mpw5_submission_0/tia_core_0/Out_2 io_analog[3] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15134 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15135 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15136 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15137 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15138 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15139 vccd1 mpw5_submission_0/eigth_mirror_0/I_In a_424970_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15140 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D117 io_analog[2] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X15141 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15142 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15143 mpw5_submission_0/outd_0/outd_stage1_0/isource_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_465060_656606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
D118 io_analog[1] vccd1 sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
X15144 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15145 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15146 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15147 mpw5_submission_1/isource_0/VM8D mpw5_submission_1/isource_0/VM9D mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X15148 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15149 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15150 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15151 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15152 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15153 mpw5_submission_0/tia_core_0/VM40D mpw5_submission_0/tia_core_0/VM39D mpw5_submission_0/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15154 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15155 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15156 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15157 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15158 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15159 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15160 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15161 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15162 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15163 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15164 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15165 mpw5_submission_1/isource_0/VM12D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM11D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X15166 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15167 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15168 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15169 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15170 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15171 mpw5_submission_1/isource_0/VM22D a_171016_648702# mpw5_submission_1/isource_0/VM3D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X15172 mpw5_submission_1/isource_0/VM22D a_171016_648702# mpw5_submission_1/isource_0/VM3D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X15173 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15174 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15175 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15176 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15177 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
D119 vssd1 io_analog[1] sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
X15178 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15179 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15180 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15181 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15182 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15183 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15184 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15185 a_203650_645683# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15186 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15187 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15188 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15189 a_434420_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15190 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15191 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15192 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15193 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15194 mpw5_submission_0/eigth_mirror_0/I_In mpw5_submission_0/isource_0/VM22D a_411216_644902# vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X15195 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15196 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15197 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15198 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15199 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15200 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15201 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15202 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15203 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15204 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15205 mpw5_submission_0/eigth_mirror_0/I_out_4 mpw5_submission_0/eigth_mirror_0/I_In a_429020_636823# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15206 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15207 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15208 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15209 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15210 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15211 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15212 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_P io_analog[0] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15213 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15214 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15215 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15216 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15217 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15218 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15219 vssd1 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM36D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15220 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15221 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15222 mpw5_submission_0/tia_core_0/VM28D io_analog[3] mpw5_submission_0/outd_0/InputSignal vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15223 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15224 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15225 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15226 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15227 io_analog[5] mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15228 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15229 io_analog[6] mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/tia_core_0/Out_2 io_analog[6] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15230 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15231 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15232 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15233 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15234 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15235 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15236 a_433070_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15237 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15238 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15239 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15240 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15241 vccd1 mpw5_submission_1/eigth_mirror_0/I_In a_191520_640623# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15242 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15243 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15244 mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/V_da1_P mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15245 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15246 vccd1 a_201520_649146# a_201720_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15247 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15248 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15249 a_435770_636823# mpw5_submission_0/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15250 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15251 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15252 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15253 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15254 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15255 mpw5_submission_0/isource_0/VM3D a_411216_644902# mpw5_submission_0/isource_0/VM22D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X15256 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15257 a_188820_640623# mpw5_submission_1/eigth_mirror_0/I_In vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15258 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15259 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15260 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15261 mpw5_submission_0/isource_0/VM12D mpw5_submission_0/isource_0/VM12G vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X15262 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15263 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15264 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15265 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15266 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15267 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15268 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15269 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15270 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15271 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15272 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15273 vccd1 mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15274 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15275 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15276 mpw5_submission_1/tia_core_0/VM28D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15277 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_224860_660406# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15278 mpw5_submission_0/tia_core_0/Out_2 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15279 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15280 vccd1 io_analog[5] vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X15281 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15282 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15283 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15284 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15285 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15286 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15287 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15288 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15289 a_224238_660400# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15290 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15291 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15292 a_443850_641883# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15293 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15294 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15295 io_analog[4] vccd1 vssd1 sky130_fd_pr__res_high_po_5p73 l=4e+06u
X15296 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15297 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15298 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15299 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15300 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15301 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15302 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15303 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15304 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15305 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15306 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15307 mpw5_submission_1/eigth_mirror_0/I_In mpw5_submission_1/isource_0/VM22D a_171016_648702# vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X15308 vccd1 mpw5_submission_0/isource_0/VM8D a_430136_648079# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X15309 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da1_N mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15310 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15311 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/V_da2_N io_analog[1] mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15312 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15313 mpw5_submission_1/outd_0/V_da2_N mpw5_submission_1/outd_0/V_da1_N mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15314 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15315 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15316 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15317 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15318 a_203370_649243# a_201520_649146# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15319 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15320 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15321 vccd1 a_201520_649146# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X15322 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15323 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15324 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15325 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15326 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15327 mpw5_submission_1/tia_core_0/Out_2 mpw5_submission_1/outd_0/InputSignal io_analog[6] io_analog[6] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15328 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15329 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15330 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15331 vccd1 a_441720_645346# a_441920_645443# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15332 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15333 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15334 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15335 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15336 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15337 vccd1 a_201520_649146# a_203650_645683# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15338 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15339 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15340 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15341 a_203370_649243# a_201520_649146# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15342 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15343 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15344 vccd1 a_201520_649146# a_203370_649243# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15345 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15346 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15347 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15348 a_224860_660406# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage1_0/isource_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15349 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15350 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15351 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15352 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15353 io_analog[6] mpw5_submission_1/outd_0/InputSignal mpw5_submission_1/tia_core_0/Out_2 io_analog[6] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15354 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15355 vssd1 mpw5_submission_1/cmirror_channel_0/TIA_I_Bias1 mpw5_submission_1/tia_core_0/VM36D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15356 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15357 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15358 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15359 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15360 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15361 io_analog[1] mpw5_submission_0/outd_0/V_da2_N mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15362 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15363 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15364 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15365 io_analog[0] mpw5_submission_0/outd_0/V_da2_P mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15366 mpw5_submission_0/outd_0/InputSignal io_analog[3] mpw5_submission_0/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15367 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15368 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15369 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15370 mpw5_submission_0/outd_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_470230_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15371 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15372 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15373 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15374 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15375 mpw5_submission_1/outd_0/InputRef mpw5_submission_1/tia_core_0/VM39D vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15376 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15377 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15378 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15379 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15380 mpw5_submission_0/tia_core_0/Out_2 mpw5_submission_0/outd_0/InputSignal io_analog[3] io_analog[3] sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15381 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15382 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15383 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15384 mpw5_submission_0/isource_0/VM11D mpw5_submission_0/isource_0/VM2D mpw5_submission_0/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X15385 mpw5_submission_1/outd_0/InputSignal io_analog[6] mpw5_submission_1/tia_core_0/VM28D vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15386 mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15387 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15388 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15389 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_230030_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15390 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15391 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15392 a_470230_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15393 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15394 mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/V_da1_P mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15395 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15396 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15397 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15398 io_analog[4] mpw5_submission_1/outd_0/V_da2_P mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15399 vccd1 a_441720_645346# a_443850_641883# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15400 mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15401 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15402 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15403 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_P io_analog[4] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15404 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15405 mpw5_submission_1/tia_core_0/VM40D mpw5_submission_1/tia_core_0/VM39D mpw5_submission_1/outd_0/InputRef vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15406 a_230030_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15407 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15408 mpw5_submission_0/tia_core_0/VM28D mpw5_submission_0/tia_core_0/Disable_TIA_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15409 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15410 vssd1 mpw5_submission_0/tia_core_0/Disable_TIA_B mpw5_submission_0/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15411 mpw5_submission_1/isource_0/VM11D mpw5_submission_1/isource_0/VM2D mpw5_submission_1/isource_0/VM12D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X15412 vssd1 mpw5_submission_1/tia_core_0/Disable_TIA_B mpw5_submission_1/tia_core_0/VM40D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15413 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15414 a_465060_656606# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15415 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15416 mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out mpw5_submission_1/outd_0/V_da2_N io_analog[5] mpw5_submission_1/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15417 vssd1 mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias a_244350_659606# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15418 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15419 a_484550_655806# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias mpw5_submission_0/outd_0/outd_stage3_0/outd_stage2_0/cmirror_out vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15420 a_244350_659606# mpw5_submission_1/cmirror_channel_0/A_Out_I_Bias vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15421 vssd1 mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias a_484550_655806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15422 a_443570_645443# a_441720_645346# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15423 a_443570_645443# a_441720_645346# mpw5_submission_0/cmirror_channel_0/A_Out_I_Bias vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u

