magic
tech sky130A
magscale 1 2
timestamp 1645701277
<< locali >>
rect 9700 11420 13840 11480
rect 11360 11400 13840 11420
rect 11460 11380 13840 11400
rect 5100 7720 5220 10860
rect 11360 9200 13840 9220
rect 9700 9140 13840 9200
rect 11460 9120 13840 9140
<< metal1 >>
rect 9600 13520 9820 13600
rect 4090 13100 4100 13340
rect 4180 13100 4190 13340
rect 4220 12620 4500 13440
rect 5360 13388 5450 13422
rect 6610 13100 6620 13340
rect 5350 12620 5360 12820
rect 5440 12620 5450 12820
rect 4220 12540 4240 12620
rect 4480 12540 4500 12620
rect 4220 12480 4500 12540
rect 5360 12478 5450 12512
rect 9600 11600 9780 13520
rect 11580 12480 11820 12640
rect 9600 11520 9820 11600
rect 9600 11340 9780 11520
rect 9600 11260 9820 11340
rect 4160 10260 5000 10720
rect 5300 10260 6160 10740
rect 6360 10260 7220 10740
rect 7420 10260 8280 10740
rect 8480 10260 9340 10740
rect 9600 9340 9780 11260
rect 11580 10220 11820 10380
rect 9600 9260 9820 9340
rect 9600 9080 9780 9260
rect 9600 9000 9820 9080
rect 4150 7820 4160 8300
rect 4480 7820 4490 8300
rect 4700 7820 5620 8300
rect 5840 7820 6700 8300
rect 6900 7820 7760 8300
rect 7960 7820 8820 8300
rect 9600 7080 9780 9000
rect 11560 7960 11800 8120
rect 9600 7000 9820 7080
<< via1 >>
rect 4100 13100 4180 13340
rect 6620 13100 6676 13340
rect 5360 12620 5440 12820
rect 4240 12540 4480 12620
rect 4160 7820 4480 8300
<< metal2 >>
rect 6760 13600 9860 13860
rect 4100 13340 4180 13350
rect 6620 13340 6700 13350
rect 4180 13100 6620 13340
rect 6676 13100 6700 13340
rect 4100 13090 4180 13100
rect 6620 13090 6700 13100
rect 5360 12820 5440 12830
rect 6760 12820 7000 13600
rect 4240 12620 4480 12630
rect 5320 12620 5360 12820
rect 5440 12620 7000 12820
rect 9600 12640 9860 13600
rect 13580 13460 13900 13700
rect 11180 13260 13900 13460
rect 4120 12540 4240 12620
rect 5360 12610 5440 12620
rect 4120 12300 4480 12540
rect 9800 12480 9860 12640
rect 4120 11960 6864 12300
rect 4120 8300 4480 11960
rect 4120 7820 4160 8300
rect 4160 7810 4480 7820
rect 9600 10380 9860 12480
rect 9800 10220 9860 10380
rect 9600 8120 9860 10220
rect 9800 7960 9860 8120
rect 9600 7720 9860 7960
rect 10060 13040 11360 13160
rect 11660 13040 12140 13160
rect 10060 12100 10220 13040
rect 12020 12680 12140 13040
rect 11800 12640 11920 12650
rect 11800 12470 11920 12480
rect 11160 12100 11300 12110
rect 10060 11980 11160 12100
rect 10060 10900 10220 11980
rect 11160 11970 11300 11980
rect 12320 12100 12460 12420
rect 12320 11970 12460 11980
rect 13580 11840 13900 13000
rect 11520 11640 13900 11840
rect 13580 11200 13900 11640
rect 11520 11000 13900 11200
rect 11120 10900 11240 10910
rect 10060 10780 11120 10900
rect 10060 8640 10220 10780
rect 11120 10770 11240 10780
rect 11660 10900 11780 10910
rect 11780 10780 12140 10900
rect 11660 10770 11780 10780
rect 12020 10420 12140 10780
rect 11800 10380 11920 10390
rect 11800 10210 11920 10220
rect 13580 9580 13900 11000
rect 11520 9380 13900 9580
rect 11040 8640 11180 8650
rect 10060 8460 11040 8640
rect 10060 7720 10220 8460
rect 11040 8450 11180 8460
rect 11760 8640 11900 8650
rect 11900 8460 12120 8640
rect 11760 8450 11900 8460
rect 12000 8160 12120 8460
rect 11800 8120 11920 8130
rect 11800 7950 11920 7960
rect 13580 6900 13900 9380
<< via2 >>
rect 9600 12480 9800 12640
rect 9600 10220 9800 10380
rect 9600 7960 9800 8120
rect 13580 13000 13900 13260
rect 11800 12480 11920 12640
rect 11160 11980 11300 12100
rect 12320 11980 12460 12100
rect 11120 10780 11240 10900
rect 11660 10780 11780 10900
rect 11800 10220 11920 10380
rect 11040 8460 11180 8640
rect 11760 8460 11900 8640
rect 11800 7960 11920 8120
<< metal3 >>
rect 9442 13260 13920 13280
rect 9442 13000 13580 13260
rect 13900 13000 13920 13260
rect 13570 12995 13910 13000
rect 9590 12640 9810 12645
rect 11790 12640 11930 12645
rect 9590 12480 9600 12640
rect 9800 12480 11800 12640
rect 11920 12480 11930 12640
rect 9590 12475 9810 12480
rect 11790 12475 11930 12480
rect 11150 12100 11310 12105
rect 12310 12100 12470 12105
rect 11150 11980 11160 12100
rect 11300 11980 12320 12100
rect 12460 11980 12470 12100
rect 11150 11975 11310 11980
rect 12310 11975 12470 11980
rect 11110 10900 11250 10905
rect 11650 10900 11790 10905
rect 11110 10780 11120 10900
rect 11240 10780 11660 10900
rect 11780 10780 11790 10900
rect 11110 10775 11250 10780
rect 11650 10775 11790 10780
rect 9590 10380 9810 10385
rect 11790 10380 11930 10385
rect 9590 10220 9600 10380
rect 9800 10220 11800 10380
rect 11920 10220 11930 10380
rect 9590 10215 9810 10220
rect 11790 10215 11930 10220
rect 11030 8640 11190 8645
rect 11750 8640 11910 8645
rect 11030 8460 11040 8640
rect 11180 8460 11760 8640
rect 11900 8460 11910 8640
rect 11030 8455 11190 8460
rect 11750 8455 11910 8460
rect 9590 8120 9810 8125
rect 11790 8120 11930 8125
rect 9590 7960 9600 8120
rect 9800 7960 11800 8120
rect 11920 7960 11930 8120
rect 9590 7955 9810 7960
rect 11790 7955 11930 7960
use isource_cmirror  isource_cmirror_0 ~/code/asic/layout/isource
timestamp 1645630008
transform 1 0 9700 0 1 11420
box 0 0 2044 2280
use isource_cmirror  isource_cmirror_1
timestamp 1645630008
transform 1 0 9700 0 1 9160
box 0 0 2044 2280
use isource_cmirror  isource_cmirror_2
timestamp 1645630008
transform 1 0 9700 0 1 6900
box 0 0 2044 2280
use isource_cmirror  isource_cmirror_3
timestamp 1645630008
transform 1 0 11740 0 1 11420
box 0 0 2044 2280
use isource_cmirror  isource_cmirror_4
timestamp 1645630008
transform 1 0 11740 0 1 9160
box 0 0 2044 2280
use isource_cmirror  isource_cmirror_5
timestamp 1645630008
transform 1 0 11740 0 1 6900
box 0 0 2044 2280
use sky130_fd_pr__nfet_01v8_WY4VMC  sky130_fd_pr__nfet_01v8_WY4VMC_2
timestamp 1645614240
transform 1 0 5405 0 1 12950
box -1425 -610 1425 610
use sky130_fd_pr__res_xhigh_po_1p41_BQY2W7  sky130_fd_pr__res_xhigh_po_1p41_BQY2W7_0
timestamp 1645462850
transform 1 0 7322 0 1 9278
box -2162 -1598 2162 1598
use sky130_fd_pr__res_xhigh_po_1p41_J2NVFM  sky130_fd_pr__res_xhigh_po_1p41_J2NVFM_0
timestamp 1645628777
transform 1 0 4592 0 1 9278
box -572 -1598 572 1598
<< end >>
