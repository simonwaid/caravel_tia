magic
tech sky130A
magscale 1 2
timestamp 1646921651
<< metal1 >>
rect 90 2440 2540 2500
rect 174 2251 184 2411
rect 236 2251 246 2411
rect 366 2251 376 2411
rect 428 2251 438 2411
rect 558 2251 568 2411
rect 620 2251 630 2411
rect 750 2251 760 2411
rect 812 2251 822 2411
rect 942 2251 952 2411
rect 1004 2251 1014 2411
rect 1134 2251 1144 2411
rect 1196 2251 1206 2411
rect 1326 2251 1336 2411
rect 1388 2251 1398 2411
rect 1518 2251 1528 2411
rect 1580 2251 1590 2411
rect 1710 2251 1720 2411
rect 1772 2251 1782 2411
rect 1902 2251 1912 2411
rect 1964 2251 1974 2411
rect 2094 2251 2104 2411
rect 2156 2251 2166 2411
rect 2286 2251 2296 2411
rect 2348 2251 2358 2411
rect 2478 2251 2488 2411
rect 2540 2251 2550 2411
rect 78 2011 88 2171
rect 140 2011 150 2171
rect 270 2011 280 2171
rect 332 2011 342 2171
rect 462 2011 472 2171
rect 524 2011 534 2171
rect 654 2011 664 2171
rect 716 2011 726 2171
rect 846 2011 856 2171
rect 908 2011 918 2171
rect 1038 2011 1048 2171
rect 1100 2011 1110 2171
rect 1230 2011 1240 2171
rect 1292 2011 1302 2171
rect 1422 2011 1432 2171
rect 1484 2011 1494 2171
rect 1614 2011 1624 2171
rect 1676 2011 1686 2171
rect 1806 2011 1816 2171
rect 1868 2011 1878 2171
rect 1998 2011 2008 2171
rect 2060 2011 2070 2171
rect 2190 2011 2200 2171
rect 2252 2011 2262 2171
rect 2382 2011 2392 2171
rect 2444 2011 2454 2171
rect 90 1830 2540 1980
rect 78 1633 88 1793
rect 140 1633 150 1793
rect 270 1633 280 1793
rect 332 1633 342 1793
rect 462 1633 472 1793
rect 524 1633 534 1793
rect 654 1633 664 1793
rect 716 1633 726 1793
rect 846 1633 856 1793
rect 908 1633 918 1793
rect 1038 1633 1048 1793
rect 1100 1633 1110 1793
rect 1230 1633 1240 1793
rect 1292 1633 1302 1793
rect 1422 1633 1432 1793
rect 1484 1633 1494 1793
rect 1614 1633 1624 1793
rect 1676 1633 1686 1793
rect 1806 1633 1816 1793
rect 1868 1633 1878 1793
rect 1998 1633 2008 1793
rect 2060 1633 2070 1793
rect 2190 1633 2200 1793
rect 2252 1633 2262 1793
rect 2382 1633 2392 1793
rect 2444 1633 2454 1793
rect 174 1393 184 1553
rect 236 1393 246 1553
rect 366 1393 376 1553
rect 428 1393 438 1553
rect 558 1393 568 1553
rect 620 1393 630 1553
rect 750 1393 760 1553
rect 812 1393 822 1553
rect 942 1393 952 1553
rect 1004 1393 1014 1553
rect 1134 1393 1144 1553
rect 1196 1393 1206 1553
rect 1326 1393 1336 1553
rect 1388 1393 1398 1553
rect 1518 1393 1528 1553
rect 1580 1393 1590 1553
rect 1710 1393 1720 1553
rect 1772 1393 1782 1553
rect 1902 1393 1912 1553
rect 1964 1393 1974 1553
rect 2094 1393 2104 1553
rect 2156 1393 2166 1553
rect 2286 1393 2296 1553
rect 2348 1393 2358 1553
rect 2478 1393 2488 1553
rect 2540 1393 2550 1553
rect 90 1210 2540 1360
rect 174 1015 184 1175
rect 236 1015 246 1175
rect 366 1015 376 1175
rect 428 1015 438 1175
rect 558 1015 568 1175
rect 620 1015 630 1175
rect 750 1015 760 1175
rect 812 1015 822 1175
rect 942 1015 952 1175
rect 1004 1015 1014 1175
rect 1134 1015 1144 1175
rect 1196 1015 1206 1175
rect 1326 1015 1336 1175
rect 1388 1015 1398 1175
rect 1518 1015 1528 1175
rect 1580 1015 1590 1175
rect 1710 1015 1720 1175
rect 1772 1015 1782 1175
rect 1902 1015 1912 1175
rect 1964 1015 1974 1175
rect 2094 1015 2104 1175
rect 2156 1015 2166 1175
rect 2286 1015 2296 1175
rect 2348 1015 2358 1175
rect 2478 1015 2488 1175
rect 2540 1015 2550 1175
rect 78 775 88 935
rect 140 775 150 935
rect 270 775 280 935
rect 332 775 342 935
rect 462 775 472 935
rect 524 775 534 935
rect 654 775 664 935
rect 716 775 726 935
rect 846 775 856 935
rect 908 775 918 935
rect 1038 775 1048 935
rect 1100 775 1110 935
rect 1230 775 1240 935
rect 1292 775 1302 935
rect 1422 775 1432 935
rect 1484 775 1494 935
rect 1614 775 1624 935
rect 1676 775 1686 935
rect 1806 775 1816 935
rect 1868 775 1878 935
rect 1998 775 2008 935
rect 2060 775 2070 935
rect 2190 775 2200 935
rect 2252 775 2262 935
rect 2382 775 2392 935
rect 2444 775 2454 935
rect 90 590 2540 740
rect 78 397 88 557
rect 140 397 150 557
rect 270 397 280 557
rect 332 397 342 557
rect 462 397 472 557
rect 524 397 534 557
rect 654 397 664 557
rect 716 397 726 557
rect 846 397 856 557
rect 908 397 918 557
rect 1038 397 1048 557
rect 1100 397 1110 557
rect 1230 397 1240 557
rect 1292 397 1302 557
rect 1422 397 1432 557
rect 1484 397 1494 557
rect 1614 397 1624 557
rect 1676 397 1686 557
rect 1806 397 1816 557
rect 1868 397 1878 557
rect 1998 397 2008 557
rect 2060 397 2070 557
rect 2190 397 2200 557
rect 2252 397 2262 557
rect 2382 397 2392 557
rect 2444 397 2454 557
rect 174 157 184 317
rect 236 157 246 317
rect 366 157 376 317
rect 428 157 438 317
rect 558 157 568 317
rect 620 157 630 317
rect 750 157 760 317
rect 812 157 822 317
rect 942 157 952 317
rect 1004 157 1014 317
rect 1134 157 1144 317
rect 1196 157 1206 317
rect 1326 157 1336 317
rect 1388 157 1398 317
rect 1518 157 1528 317
rect 1580 157 1590 317
rect 1710 157 1720 317
rect 1772 157 1782 317
rect 1902 157 1912 317
rect 1964 157 1974 317
rect 2094 157 2104 317
rect 2156 157 2166 317
rect 2286 157 2296 317
rect 2348 157 2358 317
rect 2478 157 2488 317
rect 2540 157 2550 317
rect 90 70 2540 120
<< via1 >>
rect 184 2251 236 2411
rect 376 2251 428 2411
rect 568 2251 620 2411
rect 760 2251 812 2411
rect 952 2251 1004 2411
rect 1144 2251 1196 2411
rect 1336 2251 1388 2411
rect 1528 2251 1580 2411
rect 1720 2251 1772 2411
rect 1912 2251 1964 2411
rect 2104 2251 2156 2411
rect 2296 2251 2348 2411
rect 2488 2251 2540 2411
rect 88 2011 140 2171
rect 280 2011 332 2171
rect 472 2011 524 2171
rect 664 2011 716 2171
rect 856 2011 908 2171
rect 1048 2011 1100 2171
rect 1240 2011 1292 2171
rect 1432 2011 1484 2171
rect 1624 2011 1676 2171
rect 1816 2011 1868 2171
rect 2008 2011 2060 2171
rect 2200 2011 2252 2171
rect 2392 2011 2444 2171
rect 88 1633 140 1793
rect 280 1633 332 1793
rect 472 1633 524 1793
rect 664 1633 716 1793
rect 856 1633 908 1793
rect 1048 1633 1100 1793
rect 1240 1633 1292 1793
rect 1432 1633 1484 1793
rect 1624 1633 1676 1793
rect 1816 1633 1868 1793
rect 2008 1633 2060 1793
rect 2200 1633 2252 1793
rect 2392 1633 2444 1793
rect 184 1393 236 1553
rect 376 1393 428 1553
rect 568 1393 620 1553
rect 760 1393 812 1553
rect 952 1393 1004 1553
rect 1144 1393 1196 1553
rect 1336 1393 1388 1553
rect 1528 1393 1580 1553
rect 1720 1393 1772 1553
rect 1912 1393 1964 1553
rect 2104 1393 2156 1553
rect 2296 1393 2348 1553
rect 2488 1393 2540 1553
rect 184 1015 236 1175
rect 376 1015 428 1175
rect 568 1015 620 1175
rect 760 1015 812 1175
rect 952 1015 1004 1175
rect 1144 1015 1196 1175
rect 1336 1015 1388 1175
rect 1528 1015 1580 1175
rect 1720 1015 1772 1175
rect 1912 1015 1964 1175
rect 2104 1015 2156 1175
rect 2296 1015 2348 1175
rect 2488 1015 2540 1175
rect 88 775 140 935
rect 280 775 332 935
rect 472 775 524 935
rect 664 775 716 935
rect 856 775 908 935
rect 1048 775 1100 935
rect 1240 775 1292 935
rect 1432 775 1484 935
rect 1624 775 1676 935
rect 1816 775 1868 935
rect 2008 775 2060 935
rect 2200 775 2252 935
rect 2392 775 2444 935
rect 88 397 140 557
rect 280 397 332 557
rect 472 397 524 557
rect 664 397 716 557
rect 856 397 908 557
rect 1048 397 1100 557
rect 1240 397 1292 557
rect 1432 397 1484 557
rect 1624 397 1676 557
rect 1816 397 1868 557
rect 2008 397 2060 557
rect 2200 397 2252 557
rect 2392 397 2444 557
rect 184 157 236 317
rect 376 157 428 317
rect 568 157 620 317
rect 760 157 812 317
rect 952 157 1004 317
rect 1144 157 1196 317
rect 1336 157 1388 317
rect 1528 157 1580 317
rect 1720 157 1772 317
rect 1912 157 1964 317
rect 2104 157 2156 317
rect 2296 157 2348 317
rect 2488 157 2540 317
<< metal2 >>
rect 184 2411 236 2421
rect 184 2241 236 2251
rect 376 2411 428 2421
rect 376 2241 428 2251
rect 568 2411 620 2421
rect 568 2241 620 2251
rect 760 2411 812 2421
rect 760 2241 812 2251
rect 952 2411 1004 2421
rect 952 2241 1004 2251
rect 1144 2411 1196 2421
rect 1144 2241 1196 2251
rect 1336 2411 1388 2421
rect 1336 2241 1388 2251
rect 1528 2411 1580 2421
rect 1528 2241 1580 2251
rect 1720 2411 1772 2421
rect 1720 2241 1772 2251
rect 1912 2411 1964 2421
rect 1912 2241 1964 2251
rect 2104 2411 2156 2421
rect 2104 2241 2156 2251
rect 2296 2411 2348 2421
rect 2296 2241 2348 2251
rect 2488 2411 2540 2421
rect 2488 2241 2540 2251
rect 88 2171 140 2181
rect 88 2001 140 2011
rect 280 2171 332 2181
rect 280 2001 332 2011
rect 472 2171 524 2181
rect 472 2001 524 2011
rect 664 2171 716 2181
rect 664 2001 716 2011
rect 856 2171 908 2181
rect 856 2001 908 2011
rect 1048 2171 1100 2181
rect 1048 2001 1100 2011
rect 1240 2171 1292 2181
rect 1240 2001 1292 2011
rect 1432 2171 1484 2181
rect 1432 2001 1484 2011
rect 1624 2171 1676 2181
rect 1624 2001 1676 2011
rect 1816 2171 1868 2181
rect 1816 2001 1868 2011
rect 2008 2171 2060 2181
rect 2008 2001 2060 2011
rect 2200 2171 2252 2181
rect 2200 2001 2252 2011
rect 2392 2171 2444 2181
rect 2392 2001 2444 2011
rect 88 1793 140 1803
rect 88 1623 140 1633
rect 280 1793 332 1803
rect 280 1623 332 1633
rect 472 1793 524 1803
rect 472 1623 524 1633
rect 664 1793 716 1803
rect 664 1623 716 1633
rect 856 1793 908 1803
rect 856 1623 908 1633
rect 1048 1793 1100 1803
rect 1048 1623 1100 1633
rect 1240 1793 1292 1803
rect 1240 1623 1292 1633
rect 1432 1793 1484 1803
rect 1432 1623 1484 1633
rect 1624 1793 1676 1803
rect 1624 1623 1676 1633
rect 1816 1793 1868 1803
rect 1816 1623 1868 1633
rect 2008 1793 2060 1803
rect 2008 1623 2060 1633
rect 2200 1793 2252 1803
rect 2200 1623 2252 1633
rect 2392 1793 2444 1803
rect 2392 1623 2444 1633
rect 184 1553 236 1563
rect 184 1383 236 1393
rect 376 1553 428 1563
rect 376 1383 428 1393
rect 568 1553 620 1563
rect 568 1383 620 1393
rect 760 1553 812 1563
rect 760 1383 812 1393
rect 952 1553 1004 1563
rect 952 1383 1004 1393
rect 1144 1553 1196 1563
rect 1144 1383 1196 1393
rect 1336 1553 1388 1563
rect 1336 1383 1388 1393
rect 1528 1553 1580 1563
rect 1528 1383 1580 1393
rect 1720 1553 1772 1563
rect 1720 1383 1772 1393
rect 1912 1553 1964 1563
rect 1912 1383 1964 1393
rect 2104 1553 2156 1563
rect 2104 1383 2156 1393
rect 2296 1553 2348 1563
rect 2296 1383 2348 1393
rect 2488 1553 2540 1563
rect 2488 1383 2540 1393
rect 184 1175 236 1185
rect 184 1005 236 1015
rect 376 1175 428 1185
rect 376 1005 428 1015
rect 568 1175 620 1185
rect 568 1005 620 1015
rect 760 1175 812 1185
rect 760 1005 812 1015
rect 952 1175 1004 1185
rect 952 1005 1004 1015
rect 1144 1175 1196 1185
rect 1144 1005 1196 1015
rect 1336 1175 1388 1185
rect 1336 1005 1388 1015
rect 1528 1175 1580 1185
rect 1528 1005 1580 1015
rect 1720 1175 1772 1185
rect 1720 1005 1772 1015
rect 1912 1175 1964 1185
rect 1912 1005 1964 1015
rect 2104 1175 2156 1185
rect 2104 1005 2156 1015
rect 2296 1175 2348 1185
rect 2296 1005 2348 1015
rect 2488 1175 2540 1185
rect 2488 1005 2540 1015
rect 88 935 140 945
rect 88 765 140 775
rect 280 935 332 945
rect 280 765 332 775
rect 472 935 524 945
rect 472 765 524 775
rect 664 935 716 945
rect 664 765 716 775
rect 856 935 908 945
rect 856 765 908 775
rect 1048 935 1100 945
rect 1048 765 1100 775
rect 1240 935 1292 945
rect 1240 765 1292 775
rect 1432 935 1484 945
rect 1432 765 1484 775
rect 1624 935 1676 945
rect 1624 765 1676 775
rect 1816 935 1868 945
rect 1816 765 1868 775
rect 2008 935 2060 945
rect 2008 765 2060 775
rect 2200 935 2252 945
rect 2200 765 2252 775
rect 2392 935 2444 945
rect 2392 765 2444 775
rect 88 557 140 567
rect 88 387 140 397
rect 280 557 332 567
rect 280 387 332 397
rect 472 557 524 567
rect 472 387 524 397
rect 664 557 716 567
rect 664 387 716 397
rect 856 557 908 567
rect 856 387 908 397
rect 1048 557 1100 567
rect 1048 387 1100 397
rect 1240 557 1292 567
rect 1240 387 1292 397
rect 1432 557 1484 567
rect 1432 387 1484 397
rect 1624 557 1676 567
rect 1624 387 1676 397
rect 1816 557 1868 567
rect 1816 387 1868 397
rect 2008 557 2060 567
rect 2008 387 2060 397
rect 2200 557 2252 567
rect 2200 387 2252 397
rect 2392 557 2444 567
rect 2392 387 2444 397
rect 184 317 236 327
rect 184 147 236 157
rect 376 317 428 327
rect 376 147 428 157
rect 568 317 620 327
rect 568 147 620 157
rect 760 317 812 327
rect 760 147 812 157
rect 952 317 1004 327
rect 952 147 1004 157
rect 1144 317 1196 327
rect 1144 147 1196 157
rect 1336 317 1388 327
rect 1336 147 1388 157
rect 1528 317 1580 327
rect 1528 147 1580 157
rect 1720 317 1772 327
rect 1720 147 1772 157
rect 1912 317 1964 327
rect 1912 147 1964 157
rect 2104 317 2156 327
rect 2104 147 2156 157
rect 2296 317 2348 327
rect 2296 147 2348 157
rect 2488 317 2540 327
rect 2488 147 2540 157
use sky130_fd_pr__nfet_01v8_RRWALQ  sky130_fd_pr__nfet_01v8_RRWALQ_0
timestamp 1646921651
transform 1 0 1314 0 1 1284
box -1367 -1337 1367 1337
<< end >>
