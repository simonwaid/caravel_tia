magic
tech sky130A
magscale 1 2
timestamp 1647254192
<< error_p >>
rect -1205 581 -1147 587
rect -1009 581 -951 587
rect -813 581 -755 587
rect -617 581 -559 587
rect -421 581 -363 587
rect -225 581 -167 587
rect -29 581 29 587
rect 167 581 225 587
rect 363 581 421 587
rect 559 581 617 587
rect 755 581 813 587
rect 951 581 1009 587
rect 1147 581 1205 587
rect -1205 547 -1193 581
rect -1009 547 -997 581
rect -813 547 -801 581
rect -617 547 -605 581
rect -421 547 -409 581
rect -225 547 -213 581
rect -29 547 -17 581
rect 167 547 179 581
rect 363 547 375 581
rect 559 547 571 581
rect 755 547 767 581
rect 951 547 963 581
rect 1147 547 1159 581
rect -1205 541 -1147 547
rect -1009 541 -951 547
rect -813 541 -755 547
rect -617 541 -559 547
rect -421 541 -363 547
rect -225 541 -167 547
rect -29 541 29 547
rect 167 541 225 547
rect 363 541 421 547
rect 559 541 617 547
rect 755 541 813 547
rect 951 541 1009 547
rect 1147 541 1205 547
rect -1107 71 -1049 77
rect -911 71 -853 77
rect -715 71 -657 77
rect -519 71 -461 77
rect -323 71 -265 77
rect -127 71 -69 77
rect 69 71 127 77
rect 265 71 323 77
rect 461 71 519 77
rect 657 71 715 77
rect 853 71 911 77
rect 1049 71 1107 77
rect -1107 37 -1095 71
rect -911 37 -899 71
rect -715 37 -703 71
rect -519 37 -507 71
rect -323 37 -311 71
rect -127 37 -115 71
rect 69 37 81 71
rect 265 37 277 71
rect 461 37 473 71
rect 657 37 669 71
rect 853 37 865 71
rect 1049 37 1061 71
rect -1107 31 -1049 37
rect -911 31 -853 37
rect -715 31 -657 37
rect -519 31 -461 37
rect -323 31 -265 37
rect -127 31 -69 37
rect 69 31 127 37
rect 265 31 323 37
rect 461 31 519 37
rect 657 31 715 37
rect 853 31 911 37
rect 1049 31 1107 37
rect -1107 -37 -1049 -31
rect -911 -37 -853 -31
rect -715 -37 -657 -31
rect -519 -37 -461 -31
rect -323 -37 -265 -31
rect -127 -37 -69 -31
rect 69 -37 127 -31
rect 265 -37 323 -31
rect 461 -37 519 -31
rect 657 -37 715 -31
rect 853 -37 911 -31
rect 1049 -37 1107 -31
rect -1107 -71 -1095 -37
rect -911 -71 -899 -37
rect -715 -71 -703 -37
rect -519 -71 -507 -37
rect -323 -71 -311 -37
rect -127 -71 -115 -37
rect 69 -71 81 -37
rect 265 -71 277 -37
rect 461 -71 473 -37
rect 657 -71 669 -37
rect 853 -71 865 -37
rect 1049 -71 1061 -37
rect -1107 -77 -1049 -71
rect -911 -77 -853 -71
rect -715 -77 -657 -71
rect -519 -77 -461 -71
rect -323 -77 -265 -71
rect -127 -77 -69 -71
rect 69 -77 127 -71
rect 265 -77 323 -71
rect 461 -77 519 -71
rect 657 -77 715 -71
rect 853 -77 911 -71
rect 1049 -77 1107 -71
rect -1205 -547 -1147 -541
rect -1009 -547 -951 -541
rect -813 -547 -755 -541
rect -617 -547 -559 -541
rect -421 -547 -363 -541
rect -225 -547 -167 -541
rect -29 -547 29 -541
rect 167 -547 225 -541
rect 363 -547 421 -541
rect 559 -547 617 -541
rect 755 -547 813 -541
rect 951 -547 1009 -541
rect 1147 -547 1205 -541
rect -1205 -581 -1193 -547
rect -1009 -581 -997 -547
rect -813 -581 -801 -547
rect -617 -581 -605 -547
rect -421 -581 -409 -547
rect -225 -581 -213 -547
rect -29 -581 -17 -547
rect 167 -581 179 -547
rect 363 -581 375 -547
rect 559 -581 571 -547
rect 755 -581 767 -547
rect 951 -581 963 -547
rect 1147 -581 1159 -547
rect -1205 -587 -1147 -581
rect -1009 -587 -951 -581
rect -813 -587 -755 -581
rect -617 -587 -559 -581
rect -421 -587 -363 -581
rect -225 -587 -167 -581
rect -29 -587 29 -581
rect 167 -587 225 -581
rect 363 -587 421 -581
rect 559 -587 617 -581
rect 755 -587 813 -581
rect 951 -587 1009 -581
rect 1147 -587 1205 -581
<< pwell >>
rect -1392 -719 1392 719
<< nmoslvt >>
rect -1196 109 -1156 509
rect -1098 109 -1058 509
rect -1000 109 -960 509
rect -902 109 -862 509
rect -804 109 -764 509
rect -706 109 -666 509
rect -608 109 -568 509
rect -510 109 -470 509
rect -412 109 -372 509
rect -314 109 -274 509
rect -216 109 -176 509
rect -118 109 -78 509
rect -20 109 20 509
rect 78 109 118 509
rect 176 109 216 509
rect 274 109 314 509
rect 372 109 412 509
rect 470 109 510 509
rect 568 109 608 509
rect 666 109 706 509
rect 764 109 804 509
rect 862 109 902 509
rect 960 109 1000 509
rect 1058 109 1098 509
rect 1156 109 1196 509
rect -1196 -509 -1156 -109
rect -1098 -509 -1058 -109
rect -1000 -509 -960 -109
rect -902 -509 -862 -109
rect -804 -509 -764 -109
rect -706 -509 -666 -109
rect -608 -509 -568 -109
rect -510 -509 -470 -109
rect -412 -509 -372 -109
rect -314 -509 -274 -109
rect -216 -509 -176 -109
rect -118 -509 -78 -109
rect -20 -509 20 -109
rect 78 -509 118 -109
rect 176 -509 216 -109
rect 274 -509 314 -109
rect 372 -509 412 -109
rect 470 -509 510 -109
rect 568 -509 608 -109
rect 666 -509 706 -109
rect 764 -509 804 -109
rect 862 -509 902 -109
rect 960 -509 1000 -109
rect 1058 -509 1098 -109
rect 1156 -509 1196 -109
<< ndiff >>
rect -1254 497 -1196 509
rect -1254 121 -1242 497
rect -1208 121 -1196 497
rect -1254 109 -1196 121
rect -1156 497 -1098 509
rect -1156 121 -1144 497
rect -1110 121 -1098 497
rect -1156 109 -1098 121
rect -1058 497 -1000 509
rect -1058 121 -1046 497
rect -1012 121 -1000 497
rect -1058 109 -1000 121
rect -960 497 -902 509
rect -960 121 -948 497
rect -914 121 -902 497
rect -960 109 -902 121
rect -862 497 -804 509
rect -862 121 -850 497
rect -816 121 -804 497
rect -862 109 -804 121
rect -764 497 -706 509
rect -764 121 -752 497
rect -718 121 -706 497
rect -764 109 -706 121
rect -666 497 -608 509
rect -666 121 -654 497
rect -620 121 -608 497
rect -666 109 -608 121
rect -568 497 -510 509
rect -568 121 -556 497
rect -522 121 -510 497
rect -568 109 -510 121
rect -470 497 -412 509
rect -470 121 -458 497
rect -424 121 -412 497
rect -470 109 -412 121
rect -372 497 -314 509
rect -372 121 -360 497
rect -326 121 -314 497
rect -372 109 -314 121
rect -274 497 -216 509
rect -274 121 -262 497
rect -228 121 -216 497
rect -274 109 -216 121
rect -176 497 -118 509
rect -176 121 -164 497
rect -130 121 -118 497
rect -176 109 -118 121
rect -78 497 -20 509
rect -78 121 -66 497
rect -32 121 -20 497
rect -78 109 -20 121
rect 20 497 78 509
rect 20 121 32 497
rect 66 121 78 497
rect 20 109 78 121
rect 118 497 176 509
rect 118 121 130 497
rect 164 121 176 497
rect 118 109 176 121
rect 216 497 274 509
rect 216 121 228 497
rect 262 121 274 497
rect 216 109 274 121
rect 314 497 372 509
rect 314 121 326 497
rect 360 121 372 497
rect 314 109 372 121
rect 412 497 470 509
rect 412 121 424 497
rect 458 121 470 497
rect 412 109 470 121
rect 510 497 568 509
rect 510 121 522 497
rect 556 121 568 497
rect 510 109 568 121
rect 608 497 666 509
rect 608 121 620 497
rect 654 121 666 497
rect 608 109 666 121
rect 706 497 764 509
rect 706 121 718 497
rect 752 121 764 497
rect 706 109 764 121
rect 804 497 862 509
rect 804 121 816 497
rect 850 121 862 497
rect 804 109 862 121
rect 902 497 960 509
rect 902 121 914 497
rect 948 121 960 497
rect 902 109 960 121
rect 1000 497 1058 509
rect 1000 121 1012 497
rect 1046 121 1058 497
rect 1000 109 1058 121
rect 1098 497 1156 509
rect 1098 121 1110 497
rect 1144 121 1156 497
rect 1098 109 1156 121
rect 1196 497 1254 509
rect 1196 121 1208 497
rect 1242 121 1254 497
rect 1196 109 1254 121
rect -1254 -121 -1196 -109
rect -1254 -497 -1242 -121
rect -1208 -497 -1196 -121
rect -1254 -509 -1196 -497
rect -1156 -121 -1098 -109
rect -1156 -497 -1144 -121
rect -1110 -497 -1098 -121
rect -1156 -509 -1098 -497
rect -1058 -121 -1000 -109
rect -1058 -497 -1046 -121
rect -1012 -497 -1000 -121
rect -1058 -509 -1000 -497
rect -960 -121 -902 -109
rect -960 -497 -948 -121
rect -914 -497 -902 -121
rect -960 -509 -902 -497
rect -862 -121 -804 -109
rect -862 -497 -850 -121
rect -816 -497 -804 -121
rect -862 -509 -804 -497
rect -764 -121 -706 -109
rect -764 -497 -752 -121
rect -718 -497 -706 -121
rect -764 -509 -706 -497
rect -666 -121 -608 -109
rect -666 -497 -654 -121
rect -620 -497 -608 -121
rect -666 -509 -608 -497
rect -568 -121 -510 -109
rect -568 -497 -556 -121
rect -522 -497 -510 -121
rect -568 -509 -510 -497
rect -470 -121 -412 -109
rect -470 -497 -458 -121
rect -424 -497 -412 -121
rect -470 -509 -412 -497
rect -372 -121 -314 -109
rect -372 -497 -360 -121
rect -326 -497 -314 -121
rect -372 -509 -314 -497
rect -274 -121 -216 -109
rect -274 -497 -262 -121
rect -228 -497 -216 -121
rect -274 -509 -216 -497
rect -176 -121 -118 -109
rect -176 -497 -164 -121
rect -130 -497 -118 -121
rect -176 -509 -118 -497
rect -78 -121 -20 -109
rect -78 -497 -66 -121
rect -32 -497 -20 -121
rect -78 -509 -20 -497
rect 20 -121 78 -109
rect 20 -497 32 -121
rect 66 -497 78 -121
rect 20 -509 78 -497
rect 118 -121 176 -109
rect 118 -497 130 -121
rect 164 -497 176 -121
rect 118 -509 176 -497
rect 216 -121 274 -109
rect 216 -497 228 -121
rect 262 -497 274 -121
rect 216 -509 274 -497
rect 314 -121 372 -109
rect 314 -497 326 -121
rect 360 -497 372 -121
rect 314 -509 372 -497
rect 412 -121 470 -109
rect 412 -497 424 -121
rect 458 -497 470 -121
rect 412 -509 470 -497
rect 510 -121 568 -109
rect 510 -497 522 -121
rect 556 -497 568 -121
rect 510 -509 568 -497
rect 608 -121 666 -109
rect 608 -497 620 -121
rect 654 -497 666 -121
rect 608 -509 666 -497
rect 706 -121 764 -109
rect 706 -497 718 -121
rect 752 -497 764 -121
rect 706 -509 764 -497
rect 804 -121 862 -109
rect 804 -497 816 -121
rect 850 -497 862 -121
rect 804 -509 862 -497
rect 902 -121 960 -109
rect 902 -497 914 -121
rect 948 -497 960 -121
rect 902 -509 960 -497
rect 1000 -121 1058 -109
rect 1000 -497 1012 -121
rect 1046 -497 1058 -121
rect 1000 -509 1058 -497
rect 1098 -121 1156 -109
rect 1098 -497 1110 -121
rect 1144 -497 1156 -121
rect 1098 -509 1156 -497
rect 1196 -121 1254 -109
rect 1196 -497 1208 -121
rect 1242 -497 1254 -121
rect 1196 -509 1254 -497
<< ndiffc >>
rect -1242 121 -1208 497
rect -1144 121 -1110 497
rect -1046 121 -1012 497
rect -948 121 -914 497
rect -850 121 -816 497
rect -752 121 -718 497
rect -654 121 -620 497
rect -556 121 -522 497
rect -458 121 -424 497
rect -360 121 -326 497
rect -262 121 -228 497
rect -164 121 -130 497
rect -66 121 -32 497
rect 32 121 66 497
rect 130 121 164 497
rect 228 121 262 497
rect 326 121 360 497
rect 424 121 458 497
rect 522 121 556 497
rect 620 121 654 497
rect 718 121 752 497
rect 816 121 850 497
rect 914 121 948 497
rect 1012 121 1046 497
rect 1110 121 1144 497
rect 1208 121 1242 497
rect -1242 -497 -1208 -121
rect -1144 -497 -1110 -121
rect -1046 -497 -1012 -121
rect -948 -497 -914 -121
rect -850 -497 -816 -121
rect -752 -497 -718 -121
rect -654 -497 -620 -121
rect -556 -497 -522 -121
rect -458 -497 -424 -121
rect -360 -497 -326 -121
rect -262 -497 -228 -121
rect -164 -497 -130 -121
rect -66 -497 -32 -121
rect 32 -497 66 -121
rect 130 -497 164 -121
rect 228 -497 262 -121
rect 326 -497 360 -121
rect 424 -497 458 -121
rect 522 -497 556 -121
rect 620 -497 654 -121
rect 718 -497 752 -121
rect 816 -497 850 -121
rect 914 -497 948 -121
rect 1012 -497 1046 -121
rect 1110 -497 1144 -121
rect 1208 -497 1242 -121
<< psubdiff >>
rect -1356 649 -1260 683
rect 1260 649 1356 683
rect -1356 587 -1322 649
rect 1322 587 1356 649
rect -1356 -649 -1322 -587
rect 1322 -649 1356 -587
rect -1356 -683 -1260 -649
rect 1260 -683 1356 -649
<< psubdiffcont >>
rect -1260 649 1260 683
rect -1356 -587 -1322 587
rect 1322 -587 1356 587
rect -1260 -683 1260 -649
<< poly >>
rect -1209 581 -1143 597
rect -1209 547 -1193 581
rect -1159 547 -1143 581
rect -1209 531 -1143 547
rect -1013 581 -947 597
rect -1013 547 -997 581
rect -963 547 -947 581
rect -1196 509 -1156 531
rect -1098 509 -1058 535
rect -1013 531 -947 547
rect -817 581 -751 597
rect -817 547 -801 581
rect -767 547 -751 581
rect -1000 509 -960 531
rect -902 509 -862 535
rect -817 531 -751 547
rect -621 581 -555 597
rect -621 547 -605 581
rect -571 547 -555 581
rect -804 509 -764 531
rect -706 509 -666 535
rect -621 531 -555 547
rect -425 581 -359 597
rect -425 547 -409 581
rect -375 547 -359 581
rect -608 509 -568 531
rect -510 509 -470 535
rect -425 531 -359 547
rect -229 581 -163 597
rect -229 547 -213 581
rect -179 547 -163 581
rect -412 509 -372 531
rect -314 509 -274 535
rect -229 531 -163 547
rect -33 581 33 597
rect -33 547 -17 581
rect 17 547 33 581
rect -216 509 -176 531
rect -118 509 -78 535
rect -33 531 33 547
rect 163 581 229 597
rect 163 547 179 581
rect 213 547 229 581
rect -20 509 20 531
rect 78 509 118 535
rect 163 531 229 547
rect 359 581 425 597
rect 359 547 375 581
rect 409 547 425 581
rect 176 509 216 531
rect 274 509 314 535
rect 359 531 425 547
rect 555 581 621 597
rect 555 547 571 581
rect 605 547 621 581
rect 372 509 412 531
rect 470 509 510 535
rect 555 531 621 547
rect 751 581 817 597
rect 751 547 767 581
rect 801 547 817 581
rect 568 509 608 531
rect 666 509 706 535
rect 751 531 817 547
rect 947 581 1013 597
rect 947 547 963 581
rect 997 547 1013 581
rect 764 509 804 531
rect 862 509 902 535
rect 947 531 1013 547
rect 1143 581 1209 597
rect 1143 547 1159 581
rect 1193 547 1209 581
rect 960 509 1000 531
rect 1058 509 1098 535
rect 1143 531 1209 547
rect 1156 509 1196 531
rect -1196 83 -1156 109
rect -1098 87 -1058 109
rect -1111 71 -1045 87
rect -1000 83 -960 109
rect -902 87 -862 109
rect -1111 37 -1095 71
rect -1061 37 -1045 71
rect -1111 21 -1045 37
rect -915 71 -849 87
rect -804 83 -764 109
rect -706 87 -666 109
rect -915 37 -899 71
rect -865 37 -849 71
rect -915 21 -849 37
rect -719 71 -653 87
rect -608 83 -568 109
rect -510 87 -470 109
rect -719 37 -703 71
rect -669 37 -653 71
rect -719 21 -653 37
rect -523 71 -457 87
rect -412 83 -372 109
rect -314 87 -274 109
rect -523 37 -507 71
rect -473 37 -457 71
rect -523 21 -457 37
rect -327 71 -261 87
rect -216 83 -176 109
rect -118 87 -78 109
rect -327 37 -311 71
rect -277 37 -261 71
rect -327 21 -261 37
rect -131 71 -65 87
rect -20 83 20 109
rect 78 87 118 109
rect -131 37 -115 71
rect -81 37 -65 71
rect -131 21 -65 37
rect 65 71 131 87
rect 176 83 216 109
rect 274 87 314 109
rect 65 37 81 71
rect 115 37 131 71
rect 65 21 131 37
rect 261 71 327 87
rect 372 83 412 109
rect 470 87 510 109
rect 261 37 277 71
rect 311 37 327 71
rect 261 21 327 37
rect 457 71 523 87
rect 568 83 608 109
rect 666 87 706 109
rect 457 37 473 71
rect 507 37 523 71
rect 457 21 523 37
rect 653 71 719 87
rect 764 83 804 109
rect 862 87 902 109
rect 653 37 669 71
rect 703 37 719 71
rect 653 21 719 37
rect 849 71 915 87
rect 960 83 1000 109
rect 1058 87 1098 109
rect 849 37 865 71
rect 899 37 915 71
rect 849 21 915 37
rect 1045 71 1111 87
rect 1156 83 1196 109
rect 1045 37 1061 71
rect 1095 37 1111 71
rect 1045 21 1111 37
rect -1111 -37 -1045 -21
rect -1111 -71 -1095 -37
rect -1061 -71 -1045 -37
rect -1196 -109 -1156 -83
rect -1111 -87 -1045 -71
rect -915 -37 -849 -21
rect -915 -71 -899 -37
rect -865 -71 -849 -37
rect -1098 -109 -1058 -87
rect -1000 -109 -960 -83
rect -915 -87 -849 -71
rect -719 -37 -653 -21
rect -719 -71 -703 -37
rect -669 -71 -653 -37
rect -902 -109 -862 -87
rect -804 -109 -764 -83
rect -719 -87 -653 -71
rect -523 -37 -457 -21
rect -523 -71 -507 -37
rect -473 -71 -457 -37
rect -706 -109 -666 -87
rect -608 -109 -568 -83
rect -523 -87 -457 -71
rect -327 -37 -261 -21
rect -327 -71 -311 -37
rect -277 -71 -261 -37
rect -510 -109 -470 -87
rect -412 -109 -372 -83
rect -327 -87 -261 -71
rect -131 -37 -65 -21
rect -131 -71 -115 -37
rect -81 -71 -65 -37
rect -314 -109 -274 -87
rect -216 -109 -176 -83
rect -131 -87 -65 -71
rect 65 -37 131 -21
rect 65 -71 81 -37
rect 115 -71 131 -37
rect -118 -109 -78 -87
rect -20 -109 20 -83
rect 65 -87 131 -71
rect 261 -37 327 -21
rect 261 -71 277 -37
rect 311 -71 327 -37
rect 78 -109 118 -87
rect 176 -109 216 -83
rect 261 -87 327 -71
rect 457 -37 523 -21
rect 457 -71 473 -37
rect 507 -71 523 -37
rect 274 -109 314 -87
rect 372 -109 412 -83
rect 457 -87 523 -71
rect 653 -37 719 -21
rect 653 -71 669 -37
rect 703 -71 719 -37
rect 470 -109 510 -87
rect 568 -109 608 -83
rect 653 -87 719 -71
rect 849 -37 915 -21
rect 849 -71 865 -37
rect 899 -71 915 -37
rect 666 -109 706 -87
rect 764 -109 804 -83
rect 849 -87 915 -71
rect 1045 -37 1111 -21
rect 1045 -71 1061 -37
rect 1095 -71 1111 -37
rect 862 -109 902 -87
rect 960 -109 1000 -83
rect 1045 -87 1111 -71
rect 1058 -109 1098 -87
rect 1156 -109 1196 -83
rect -1196 -531 -1156 -509
rect -1209 -547 -1143 -531
rect -1098 -535 -1058 -509
rect -1000 -531 -960 -509
rect -1209 -581 -1193 -547
rect -1159 -581 -1143 -547
rect -1209 -597 -1143 -581
rect -1013 -547 -947 -531
rect -902 -535 -862 -509
rect -804 -531 -764 -509
rect -1013 -581 -997 -547
rect -963 -581 -947 -547
rect -1013 -597 -947 -581
rect -817 -547 -751 -531
rect -706 -535 -666 -509
rect -608 -531 -568 -509
rect -817 -581 -801 -547
rect -767 -581 -751 -547
rect -817 -597 -751 -581
rect -621 -547 -555 -531
rect -510 -535 -470 -509
rect -412 -531 -372 -509
rect -621 -581 -605 -547
rect -571 -581 -555 -547
rect -621 -597 -555 -581
rect -425 -547 -359 -531
rect -314 -535 -274 -509
rect -216 -531 -176 -509
rect -425 -581 -409 -547
rect -375 -581 -359 -547
rect -425 -597 -359 -581
rect -229 -547 -163 -531
rect -118 -535 -78 -509
rect -20 -531 20 -509
rect -229 -581 -213 -547
rect -179 -581 -163 -547
rect -229 -597 -163 -581
rect -33 -547 33 -531
rect 78 -535 118 -509
rect 176 -531 216 -509
rect -33 -581 -17 -547
rect 17 -581 33 -547
rect -33 -597 33 -581
rect 163 -547 229 -531
rect 274 -535 314 -509
rect 372 -531 412 -509
rect 163 -581 179 -547
rect 213 -581 229 -547
rect 163 -597 229 -581
rect 359 -547 425 -531
rect 470 -535 510 -509
rect 568 -531 608 -509
rect 359 -581 375 -547
rect 409 -581 425 -547
rect 359 -597 425 -581
rect 555 -547 621 -531
rect 666 -535 706 -509
rect 764 -531 804 -509
rect 555 -581 571 -547
rect 605 -581 621 -547
rect 555 -597 621 -581
rect 751 -547 817 -531
rect 862 -535 902 -509
rect 960 -531 1000 -509
rect 751 -581 767 -547
rect 801 -581 817 -547
rect 751 -597 817 -581
rect 947 -547 1013 -531
rect 1058 -535 1098 -509
rect 1156 -531 1196 -509
rect 947 -581 963 -547
rect 997 -581 1013 -547
rect 947 -597 1013 -581
rect 1143 -547 1209 -531
rect 1143 -581 1159 -547
rect 1193 -581 1209 -547
rect 1143 -597 1209 -581
<< polycont >>
rect -1193 547 -1159 581
rect -997 547 -963 581
rect -801 547 -767 581
rect -605 547 -571 581
rect -409 547 -375 581
rect -213 547 -179 581
rect -17 547 17 581
rect 179 547 213 581
rect 375 547 409 581
rect 571 547 605 581
rect 767 547 801 581
rect 963 547 997 581
rect 1159 547 1193 581
rect -1095 37 -1061 71
rect -899 37 -865 71
rect -703 37 -669 71
rect -507 37 -473 71
rect -311 37 -277 71
rect -115 37 -81 71
rect 81 37 115 71
rect 277 37 311 71
rect 473 37 507 71
rect 669 37 703 71
rect 865 37 899 71
rect 1061 37 1095 71
rect -1095 -71 -1061 -37
rect -899 -71 -865 -37
rect -703 -71 -669 -37
rect -507 -71 -473 -37
rect -311 -71 -277 -37
rect -115 -71 -81 -37
rect 81 -71 115 -37
rect 277 -71 311 -37
rect 473 -71 507 -37
rect 669 -71 703 -37
rect 865 -71 899 -37
rect 1061 -71 1095 -37
rect -1193 -581 -1159 -547
rect -997 -581 -963 -547
rect -801 -581 -767 -547
rect -605 -581 -571 -547
rect -409 -581 -375 -547
rect -213 -581 -179 -547
rect -17 -581 17 -547
rect 179 -581 213 -547
rect 375 -581 409 -547
rect 571 -581 605 -547
rect 767 -581 801 -547
rect 963 -581 997 -547
rect 1159 -581 1193 -547
<< locali >>
rect -1356 649 -1260 683
rect 1260 649 1356 683
rect -1356 587 -1322 649
rect 1322 587 1356 649
rect -1209 547 -1193 581
rect -1159 547 -1143 581
rect -1013 547 -997 581
rect -963 547 -947 581
rect -817 547 -801 581
rect -767 547 -751 581
rect -621 547 -605 581
rect -571 547 -555 581
rect -425 547 -409 581
rect -375 547 -359 581
rect -229 547 -213 581
rect -179 547 -163 581
rect -33 547 -17 581
rect 17 547 33 581
rect 163 547 179 581
rect 213 547 229 581
rect 359 547 375 581
rect 409 547 425 581
rect 555 547 571 581
rect 605 547 621 581
rect 751 547 767 581
rect 801 547 817 581
rect 947 547 963 581
rect 997 547 1013 581
rect 1143 547 1159 581
rect 1193 547 1209 581
rect -1242 497 -1208 513
rect -1242 105 -1208 121
rect -1144 497 -1110 513
rect -1144 105 -1110 121
rect -1046 497 -1012 513
rect -1046 105 -1012 121
rect -948 497 -914 513
rect -948 105 -914 121
rect -850 497 -816 513
rect -850 105 -816 121
rect -752 497 -718 513
rect -752 105 -718 121
rect -654 497 -620 513
rect -654 105 -620 121
rect -556 497 -522 513
rect -556 105 -522 121
rect -458 497 -424 513
rect -458 105 -424 121
rect -360 497 -326 513
rect -360 105 -326 121
rect -262 497 -228 513
rect -262 105 -228 121
rect -164 497 -130 513
rect -164 105 -130 121
rect -66 497 -32 513
rect -66 105 -32 121
rect 32 497 66 513
rect 32 105 66 121
rect 130 497 164 513
rect 130 105 164 121
rect 228 497 262 513
rect 228 105 262 121
rect 326 497 360 513
rect 326 105 360 121
rect 424 497 458 513
rect 424 105 458 121
rect 522 497 556 513
rect 522 105 556 121
rect 620 497 654 513
rect 620 105 654 121
rect 718 497 752 513
rect 718 105 752 121
rect 816 497 850 513
rect 816 105 850 121
rect 914 497 948 513
rect 914 105 948 121
rect 1012 497 1046 513
rect 1012 105 1046 121
rect 1110 497 1144 513
rect 1110 105 1144 121
rect 1208 497 1242 513
rect 1208 105 1242 121
rect -1111 37 -1095 71
rect -1061 37 -1045 71
rect -915 37 -899 71
rect -865 37 -849 71
rect -719 37 -703 71
rect -669 37 -653 71
rect -523 37 -507 71
rect -473 37 -457 71
rect -327 37 -311 71
rect -277 37 -261 71
rect -131 37 -115 71
rect -81 37 -65 71
rect 65 37 81 71
rect 115 37 131 71
rect 261 37 277 71
rect 311 37 327 71
rect 457 37 473 71
rect 507 37 523 71
rect 653 37 669 71
rect 703 37 719 71
rect 849 37 865 71
rect 899 37 915 71
rect 1045 37 1061 71
rect 1095 37 1111 71
rect -1111 -71 -1095 -37
rect -1061 -71 -1045 -37
rect -915 -71 -899 -37
rect -865 -71 -849 -37
rect -719 -71 -703 -37
rect -669 -71 -653 -37
rect -523 -71 -507 -37
rect -473 -71 -457 -37
rect -327 -71 -311 -37
rect -277 -71 -261 -37
rect -131 -71 -115 -37
rect -81 -71 -65 -37
rect 65 -71 81 -37
rect 115 -71 131 -37
rect 261 -71 277 -37
rect 311 -71 327 -37
rect 457 -71 473 -37
rect 507 -71 523 -37
rect 653 -71 669 -37
rect 703 -71 719 -37
rect 849 -71 865 -37
rect 899 -71 915 -37
rect 1045 -71 1061 -37
rect 1095 -71 1111 -37
rect -1242 -121 -1208 -105
rect -1242 -513 -1208 -497
rect -1144 -121 -1110 -105
rect -1144 -513 -1110 -497
rect -1046 -121 -1012 -105
rect -1046 -513 -1012 -497
rect -948 -121 -914 -105
rect -948 -513 -914 -497
rect -850 -121 -816 -105
rect -850 -513 -816 -497
rect -752 -121 -718 -105
rect -752 -513 -718 -497
rect -654 -121 -620 -105
rect -654 -513 -620 -497
rect -556 -121 -522 -105
rect -556 -513 -522 -497
rect -458 -121 -424 -105
rect -458 -513 -424 -497
rect -360 -121 -326 -105
rect -360 -513 -326 -497
rect -262 -121 -228 -105
rect -262 -513 -228 -497
rect -164 -121 -130 -105
rect -164 -513 -130 -497
rect -66 -121 -32 -105
rect -66 -513 -32 -497
rect 32 -121 66 -105
rect 32 -513 66 -497
rect 130 -121 164 -105
rect 130 -513 164 -497
rect 228 -121 262 -105
rect 228 -513 262 -497
rect 326 -121 360 -105
rect 326 -513 360 -497
rect 424 -121 458 -105
rect 424 -513 458 -497
rect 522 -121 556 -105
rect 522 -513 556 -497
rect 620 -121 654 -105
rect 620 -513 654 -497
rect 718 -121 752 -105
rect 718 -513 752 -497
rect 816 -121 850 -105
rect 816 -513 850 -497
rect 914 -121 948 -105
rect 914 -513 948 -497
rect 1012 -121 1046 -105
rect 1012 -513 1046 -497
rect 1110 -121 1144 -105
rect 1110 -513 1144 -497
rect 1208 -121 1242 -105
rect 1208 -513 1242 -497
rect -1209 -581 -1193 -547
rect -1159 -581 -1143 -547
rect -1013 -581 -997 -547
rect -963 -581 -947 -547
rect -817 -581 -801 -547
rect -767 -581 -751 -547
rect -621 -581 -605 -547
rect -571 -581 -555 -547
rect -425 -581 -409 -547
rect -375 -581 -359 -547
rect -229 -581 -213 -547
rect -179 -581 -163 -547
rect -33 -581 -17 -547
rect 17 -581 33 -547
rect 163 -581 179 -547
rect 213 -581 229 -547
rect 359 -581 375 -547
rect 409 -581 425 -547
rect 555 -581 571 -547
rect 605 -581 621 -547
rect 751 -581 767 -547
rect 801 -581 817 -547
rect 947 -581 963 -547
rect 997 -581 1013 -547
rect 1143 -581 1159 -547
rect 1193 -581 1209 -547
rect -1356 -649 -1322 -587
rect 1322 -649 1356 -587
rect -1356 -683 -1260 -649
rect 1260 -683 1356 -649
<< viali >>
rect -1193 547 -1159 581
rect -997 547 -963 581
rect -801 547 -767 581
rect -605 547 -571 581
rect -409 547 -375 581
rect -213 547 -179 581
rect -17 547 17 581
rect 179 547 213 581
rect 375 547 409 581
rect 571 547 605 581
rect 767 547 801 581
rect 963 547 997 581
rect 1159 547 1193 581
rect -1242 121 -1208 497
rect -1144 121 -1110 497
rect -1046 121 -1012 497
rect -948 121 -914 497
rect -850 121 -816 497
rect -752 121 -718 497
rect -654 121 -620 497
rect -556 121 -522 497
rect -458 121 -424 497
rect -360 121 -326 497
rect -262 121 -228 497
rect -164 121 -130 497
rect -66 121 -32 497
rect 32 121 66 497
rect 130 121 164 497
rect 228 121 262 497
rect 326 121 360 497
rect 424 121 458 497
rect 522 121 556 497
rect 620 121 654 497
rect 718 121 752 497
rect 816 121 850 497
rect 914 121 948 497
rect 1012 121 1046 497
rect 1110 121 1144 497
rect 1208 121 1242 497
rect -1095 37 -1061 71
rect -899 37 -865 71
rect -703 37 -669 71
rect -507 37 -473 71
rect -311 37 -277 71
rect -115 37 -81 71
rect 81 37 115 71
rect 277 37 311 71
rect 473 37 507 71
rect 669 37 703 71
rect 865 37 899 71
rect 1061 37 1095 71
rect -1095 -71 -1061 -37
rect -899 -71 -865 -37
rect -703 -71 -669 -37
rect -507 -71 -473 -37
rect -311 -71 -277 -37
rect -115 -71 -81 -37
rect 81 -71 115 -37
rect 277 -71 311 -37
rect 473 -71 507 -37
rect 669 -71 703 -37
rect 865 -71 899 -37
rect 1061 -71 1095 -37
rect -1242 -497 -1208 -121
rect -1144 -497 -1110 -121
rect -1046 -497 -1012 -121
rect -948 -497 -914 -121
rect -850 -497 -816 -121
rect -752 -497 -718 -121
rect -654 -497 -620 -121
rect -556 -497 -522 -121
rect -458 -497 -424 -121
rect -360 -497 -326 -121
rect -262 -497 -228 -121
rect -164 -497 -130 -121
rect -66 -497 -32 -121
rect 32 -497 66 -121
rect 130 -497 164 -121
rect 228 -497 262 -121
rect 326 -497 360 -121
rect 424 -497 458 -121
rect 522 -497 556 -121
rect 620 -497 654 -121
rect 718 -497 752 -121
rect 816 -497 850 -121
rect 914 -497 948 -121
rect 1012 -497 1046 -121
rect 1110 -497 1144 -121
rect 1208 -497 1242 -121
rect -1193 -581 -1159 -547
rect -997 -581 -963 -547
rect -801 -581 -767 -547
rect -605 -581 -571 -547
rect -409 -581 -375 -547
rect -213 -581 -179 -547
rect -17 -581 17 -547
rect 179 -581 213 -547
rect 375 -581 409 -547
rect 571 -581 605 -547
rect 767 -581 801 -547
rect 963 -581 997 -547
rect 1159 -581 1193 -547
<< metal1 >>
rect -1205 581 -1147 587
rect -1205 547 -1193 581
rect -1159 547 -1147 581
rect -1205 541 -1147 547
rect -1009 581 -951 587
rect -1009 547 -997 581
rect -963 547 -951 581
rect -1009 541 -951 547
rect -813 581 -755 587
rect -813 547 -801 581
rect -767 547 -755 581
rect -813 541 -755 547
rect -617 581 -559 587
rect -617 547 -605 581
rect -571 547 -559 581
rect -617 541 -559 547
rect -421 581 -363 587
rect -421 547 -409 581
rect -375 547 -363 581
rect -421 541 -363 547
rect -225 581 -167 587
rect -225 547 -213 581
rect -179 547 -167 581
rect -225 541 -167 547
rect -29 581 29 587
rect -29 547 -17 581
rect 17 547 29 581
rect -29 541 29 547
rect 167 581 225 587
rect 167 547 179 581
rect 213 547 225 581
rect 167 541 225 547
rect 363 581 421 587
rect 363 547 375 581
rect 409 547 421 581
rect 363 541 421 547
rect 559 581 617 587
rect 559 547 571 581
rect 605 547 617 581
rect 559 541 617 547
rect 755 581 813 587
rect 755 547 767 581
rect 801 547 813 581
rect 755 541 813 547
rect 951 581 1009 587
rect 951 547 963 581
rect 997 547 1009 581
rect 951 541 1009 547
rect 1147 581 1205 587
rect 1147 547 1159 581
rect 1193 547 1205 581
rect 1147 541 1205 547
rect -1248 497 -1202 509
rect -1248 121 -1242 497
rect -1208 121 -1202 497
rect -1248 109 -1202 121
rect -1150 497 -1104 509
rect -1150 121 -1144 497
rect -1110 121 -1104 497
rect -1150 109 -1104 121
rect -1052 497 -1006 509
rect -1052 121 -1046 497
rect -1012 121 -1006 497
rect -1052 109 -1006 121
rect -954 497 -908 509
rect -954 121 -948 497
rect -914 121 -908 497
rect -954 109 -908 121
rect -856 497 -810 509
rect -856 121 -850 497
rect -816 121 -810 497
rect -856 109 -810 121
rect -758 497 -712 509
rect -758 121 -752 497
rect -718 121 -712 497
rect -758 109 -712 121
rect -660 497 -614 509
rect -660 121 -654 497
rect -620 121 -614 497
rect -660 109 -614 121
rect -562 497 -516 509
rect -562 121 -556 497
rect -522 121 -516 497
rect -562 109 -516 121
rect -464 497 -418 509
rect -464 121 -458 497
rect -424 121 -418 497
rect -464 109 -418 121
rect -366 497 -320 509
rect -366 121 -360 497
rect -326 121 -320 497
rect -366 109 -320 121
rect -268 497 -222 509
rect -268 121 -262 497
rect -228 121 -222 497
rect -268 109 -222 121
rect -170 497 -124 509
rect -170 121 -164 497
rect -130 121 -124 497
rect -170 109 -124 121
rect -72 497 -26 509
rect -72 121 -66 497
rect -32 121 -26 497
rect -72 109 -26 121
rect 26 497 72 509
rect 26 121 32 497
rect 66 121 72 497
rect 26 109 72 121
rect 124 497 170 509
rect 124 121 130 497
rect 164 121 170 497
rect 124 109 170 121
rect 222 497 268 509
rect 222 121 228 497
rect 262 121 268 497
rect 222 109 268 121
rect 320 497 366 509
rect 320 121 326 497
rect 360 121 366 497
rect 320 109 366 121
rect 418 497 464 509
rect 418 121 424 497
rect 458 121 464 497
rect 418 109 464 121
rect 516 497 562 509
rect 516 121 522 497
rect 556 121 562 497
rect 516 109 562 121
rect 614 497 660 509
rect 614 121 620 497
rect 654 121 660 497
rect 614 109 660 121
rect 712 497 758 509
rect 712 121 718 497
rect 752 121 758 497
rect 712 109 758 121
rect 810 497 856 509
rect 810 121 816 497
rect 850 121 856 497
rect 810 109 856 121
rect 908 497 954 509
rect 908 121 914 497
rect 948 121 954 497
rect 908 109 954 121
rect 1006 497 1052 509
rect 1006 121 1012 497
rect 1046 121 1052 497
rect 1006 109 1052 121
rect 1104 497 1150 509
rect 1104 121 1110 497
rect 1144 121 1150 497
rect 1104 109 1150 121
rect 1202 497 1248 509
rect 1202 121 1208 497
rect 1242 121 1248 497
rect 1202 109 1248 121
rect -1107 71 -1049 77
rect -1107 37 -1095 71
rect -1061 37 -1049 71
rect -1107 31 -1049 37
rect -911 71 -853 77
rect -911 37 -899 71
rect -865 37 -853 71
rect -911 31 -853 37
rect -715 71 -657 77
rect -715 37 -703 71
rect -669 37 -657 71
rect -715 31 -657 37
rect -519 71 -461 77
rect -519 37 -507 71
rect -473 37 -461 71
rect -519 31 -461 37
rect -323 71 -265 77
rect -323 37 -311 71
rect -277 37 -265 71
rect -323 31 -265 37
rect -127 71 -69 77
rect -127 37 -115 71
rect -81 37 -69 71
rect -127 31 -69 37
rect 69 71 127 77
rect 69 37 81 71
rect 115 37 127 71
rect 69 31 127 37
rect 265 71 323 77
rect 265 37 277 71
rect 311 37 323 71
rect 265 31 323 37
rect 461 71 519 77
rect 461 37 473 71
rect 507 37 519 71
rect 461 31 519 37
rect 657 71 715 77
rect 657 37 669 71
rect 703 37 715 71
rect 657 31 715 37
rect 853 71 911 77
rect 853 37 865 71
rect 899 37 911 71
rect 853 31 911 37
rect 1049 71 1107 77
rect 1049 37 1061 71
rect 1095 37 1107 71
rect 1049 31 1107 37
rect -1107 -37 -1049 -31
rect -1107 -71 -1095 -37
rect -1061 -71 -1049 -37
rect -1107 -77 -1049 -71
rect -911 -37 -853 -31
rect -911 -71 -899 -37
rect -865 -71 -853 -37
rect -911 -77 -853 -71
rect -715 -37 -657 -31
rect -715 -71 -703 -37
rect -669 -71 -657 -37
rect -715 -77 -657 -71
rect -519 -37 -461 -31
rect -519 -71 -507 -37
rect -473 -71 -461 -37
rect -519 -77 -461 -71
rect -323 -37 -265 -31
rect -323 -71 -311 -37
rect -277 -71 -265 -37
rect -323 -77 -265 -71
rect -127 -37 -69 -31
rect -127 -71 -115 -37
rect -81 -71 -69 -37
rect -127 -77 -69 -71
rect 69 -37 127 -31
rect 69 -71 81 -37
rect 115 -71 127 -37
rect 69 -77 127 -71
rect 265 -37 323 -31
rect 265 -71 277 -37
rect 311 -71 323 -37
rect 265 -77 323 -71
rect 461 -37 519 -31
rect 461 -71 473 -37
rect 507 -71 519 -37
rect 461 -77 519 -71
rect 657 -37 715 -31
rect 657 -71 669 -37
rect 703 -71 715 -37
rect 657 -77 715 -71
rect 853 -37 911 -31
rect 853 -71 865 -37
rect 899 -71 911 -37
rect 853 -77 911 -71
rect 1049 -37 1107 -31
rect 1049 -71 1061 -37
rect 1095 -71 1107 -37
rect 1049 -77 1107 -71
rect -1248 -121 -1202 -109
rect -1248 -497 -1242 -121
rect -1208 -497 -1202 -121
rect -1248 -509 -1202 -497
rect -1150 -121 -1104 -109
rect -1150 -497 -1144 -121
rect -1110 -497 -1104 -121
rect -1150 -509 -1104 -497
rect -1052 -121 -1006 -109
rect -1052 -497 -1046 -121
rect -1012 -497 -1006 -121
rect -1052 -509 -1006 -497
rect -954 -121 -908 -109
rect -954 -497 -948 -121
rect -914 -497 -908 -121
rect -954 -509 -908 -497
rect -856 -121 -810 -109
rect -856 -497 -850 -121
rect -816 -497 -810 -121
rect -856 -509 -810 -497
rect -758 -121 -712 -109
rect -758 -497 -752 -121
rect -718 -497 -712 -121
rect -758 -509 -712 -497
rect -660 -121 -614 -109
rect -660 -497 -654 -121
rect -620 -497 -614 -121
rect -660 -509 -614 -497
rect -562 -121 -516 -109
rect -562 -497 -556 -121
rect -522 -497 -516 -121
rect -562 -509 -516 -497
rect -464 -121 -418 -109
rect -464 -497 -458 -121
rect -424 -497 -418 -121
rect -464 -509 -418 -497
rect -366 -121 -320 -109
rect -366 -497 -360 -121
rect -326 -497 -320 -121
rect -366 -509 -320 -497
rect -268 -121 -222 -109
rect -268 -497 -262 -121
rect -228 -497 -222 -121
rect -268 -509 -222 -497
rect -170 -121 -124 -109
rect -170 -497 -164 -121
rect -130 -497 -124 -121
rect -170 -509 -124 -497
rect -72 -121 -26 -109
rect -72 -497 -66 -121
rect -32 -497 -26 -121
rect -72 -509 -26 -497
rect 26 -121 72 -109
rect 26 -497 32 -121
rect 66 -497 72 -121
rect 26 -509 72 -497
rect 124 -121 170 -109
rect 124 -497 130 -121
rect 164 -497 170 -121
rect 124 -509 170 -497
rect 222 -121 268 -109
rect 222 -497 228 -121
rect 262 -497 268 -121
rect 222 -509 268 -497
rect 320 -121 366 -109
rect 320 -497 326 -121
rect 360 -497 366 -121
rect 320 -509 366 -497
rect 418 -121 464 -109
rect 418 -497 424 -121
rect 458 -497 464 -121
rect 418 -509 464 -497
rect 516 -121 562 -109
rect 516 -497 522 -121
rect 556 -497 562 -121
rect 516 -509 562 -497
rect 614 -121 660 -109
rect 614 -497 620 -121
rect 654 -497 660 -121
rect 614 -509 660 -497
rect 712 -121 758 -109
rect 712 -497 718 -121
rect 752 -497 758 -121
rect 712 -509 758 -497
rect 810 -121 856 -109
rect 810 -497 816 -121
rect 850 -497 856 -121
rect 810 -509 856 -497
rect 908 -121 954 -109
rect 908 -497 914 -121
rect 948 -497 954 -121
rect 908 -509 954 -497
rect 1006 -121 1052 -109
rect 1006 -497 1012 -121
rect 1046 -497 1052 -121
rect 1006 -509 1052 -497
rect 1104 -121 1150 -109
rect 1104 -497 1110 -121
rect 1144 -497 1150 -121
rect 1104 -509 1150 -497
rect 1202 -121 1248 -109
rect 1202 -497 1208 -121
rect 1242 -497 1248 -121
rect 1202 -509 1248 -497
rect -1205 -547 -1147 -541
rect -1205 -581 -1193 -547
rect -1159 -581 -1147 -547
rect -1205 -587 -1147 -581
rect -1009 -547 -951 -541
rect -1009 -581 -997 -547
rect -963 -581 -951 -547
rect -1009 -587 -951 -581
rect -813 -547 -755 -541
rect -813 -581 -801 -547
rect -767 -581 -755 -547
rect -813 -587 -755 -581
rect -617 -547 -559 -541
rect -617 -581 -605 -547
rect -571 -581 -559 -547
rect -617 -587 -559 -581
rect -421 -547 -363 -541
rect -421 -581 -409 -547
rect -375 -581 -363 -547
rect -421 -587 -363 -581
rect -225 -547 -167 -541
rect -225 -581 -213 -547
rect -179 -581 -167 -547
rect -225 -587 -167 -581
rect -29 -547 29 -541
rect -29 -581 -17 -547
rect 17 -581 29 -547
rect -29 -587 29 -581
rect 167 -547 225 -541
rect 167 -581 179 -547
rect 213 -581 225 -547
rect 167 -587 225 -581
rect 363 -547 421 -541
rect 363 -581 375 -547
rect 409 -581 421 -547
rect 363 -587 421 -581
rect 559 -547 617 -541
rect 559 -581 571 -547
rect 605 -581 617 -547
rect 559 -587 617 -581
rect 755 -547 813 -541
rect 755 -581 767 -547
rect 801 -581 813 -547
rect 755 -587 813 -581
rect 951 -547 1009 -541
rect 951 -581 963 -547
rect 997 -581 1009 -547
rect 951 -587 1009 -581
rect 1147 -547 1205 -541
rect 1147 -581 1159 -547
rect 1193 -581 1205 -547
rect 1147 -587 1205 -581
<< properties >>
string FIXED_BBOX -1339 -666 1339 666
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 0.2 m 2 nf 25 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
