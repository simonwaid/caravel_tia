magic
tech sky130A
timestamp 1646921651
<< pwell >>
rect -1816 -169 1816 169
<< psubdiff >>
rect -1798 134 -1750 151
rect -1544 134 -1496 151
rect -1798 103 -1781 134
rect -1513 103 -1496 134
rect -1798 -134 -1781 -103
rect -1513 -134 -1496 -103
rect -1798 -151 -1750 -134
rect -1544 -151 -1496 -134
rect -1432 134 -1384 151
rect -1178 134 -1130 151
rect -1432 103 -1415 134
rect -1147 103 -1130 134
rect -1432 -134 -1415 -103
rect -1147 -134 -1130 -103
rect -1432 -151 -1384 -134
rect -1178 -151 -1130 -134
rect -1066 134 -1018 151
rect -812 134 -764 151
rect -1066 103 -1049 134
rect -781 103 -764 134
rect -1066 -134 -1049 -103
rect -781 -134 -764 -103
rect -1066 -151 -1018 -134
rect -812 -151 -764 -134
rect -700 134 -652 151
rect -446 134 -398 151
rect -700 103 -683 134
rect -415 103 -398 134
rect -700 -134 -683 -103
rect -415 -134 -398 -103
rect -700 -151 -652 -134
rect -446 -151 -398 -134
rect -334 134 -286 151
rect -80 134 -32 151
rect -334 103 -317 134
rect -49 103 -32 134
rect -334 -134 -317 -103
rect -49 -134 -32 -103
rect -334 -151 -286 -134
rect -80 -151 -32 -134
rect 32 134 80 151
rect 286 134 334 151
rect 32 103 49 134
rect 317 103 334 134
rect 32 -134 49 -103
rect 317 -134 334 -103
rect 32 -151 80 -134
rect 286 -151 334 -134
rect 398 134 446 151
rect 652 134 700 151
rect 398 103 415 134
rect 683 103 700 134
rect 398 -134 415 -103
rect 683 -134 700 -103
rect 398 -151 446 -134
rect 652 -151 700 -134
rect 764 134 812 151
rect 1018 134 1066 151
rect 764 103 781 134
rect 1049 103 1066 134
rect 764 -134 781 -103
rect 1049 -134 1066 -103
rect 764 -151 812 -134
rect 1018 -151 1066 -134
rect 1130 134 1178 151
rect 1384 134 1432 151
rect 1130 103 1147 134
rect 1415 103 1432 134
rect 1130 -134 1147 -103
rect 1415 -134 1432 -103
rect 1130 -151 1178 -134
rect 1384 -151 1432 -134
rect 1496 134 1544 151
rect 1750 134 1798 151
rect 1496 103 1513 134
rect 1781 103 1798 134
rect 1496 -134 1513 -103
rect 1781 -134 1798 -103
rect 1496 -151 1544 -134
rect 1750 -151 1798 -134
<< psubdiffcont >>
rect -1750 134 -1544 151
rect -1798 -103 -1781 103
rect -1513 -103 -1496 103
rect -1750 -151 -1544 -134
rect -1384 134 -1178 151
rect -1432 -103 -1415 103
rect -1147 -103 -1130 103
rect -1384 -151 -1178 -134
rect -1018 134 -812 151
rect -1066 -103 -1049 103
rect -781 -103 -764 103
rect -1018 -151 -812 -134
rect -652 134 -446 151
rect -700 -103 -683 103
rect -415 -103 -398 103
rect -652 -151 -446 -134
rect -286 134 -80 151
rect -334 -103 -317 103
rect -49 -103 -32 103
rect -286 -151 -80 -134
rect 80 134 286 151
rect 32 -103 49 103
rect 317 -103 334 103
rect 80 -151 286 -134
rect 446 134 652 151
rect 398 -103 415 103
rect 683 -103 700 103
rect 446 -151 652 -134
rect 812 134 1018 151
rect 764 -103 781 103
rect 1049 -103 1066 103
rect 812 -151 1018 -134
rect 1178 134 1384 151
rect 1130 -103 1147 103
rect 1415 -103 1432 103
rect 1178 -151 1384 -134
rect 1544 134 1750 151
rect 1496 -103 1513 103
rect 1781 -103 1798 103
rect 1544 -151 1750 -134
<< ndiode >>
rect -1747 94 -1547 100
rect -1747 -94 -1741 94
rect -1553 -94 -1547 94
rect -1747 -100 -1547 -94
rect -1381 94 -1181 100
rect -1381 -94 -1375 94
rect -1187 -94 -1181 94
rect -1381 -100 -1181 -94
rect -1015 94 -815 100
rect -1015 -94 -1009 94
rect -821 -94 -815 94
rect -1015 -100 -815 -94
rect -649 94 -449 100
rect -649 -94 -643 94
rect -455 -94 -449 94
rect -649 -100 -449 -94
rect -283 94 -83 100
rect -283 -94 -277 94
rect -89 -94 -83 94
rect -283 -100 -83 -94
rect 83 94 283 100
rect 83 -94 89 94
rect 277 -94 283 94
rect 83 -100 283 -94
rect 449 94 649 100
rect 449 -94 455 94
rect 643 -94 649 94
rect 449 -100 649 -94
rect 815 94 1015 100
rect 815 -94 821 94
rect 1009 -94 1015 94
rect 815 -100 1015 -94
rect 1181 94 1381 100
rect 1181 -94 1187 94
rect 1375 -94 1381 94
rect 1181 -100 1381 -94
rect 1547 94 1747 100
rect 1547 -94 1553 94
rect 1741 -94 1747 94
rect 1547 -100 1747 -94
<< ndiodec >>
rect -1741 -94 -1553 94
rect -1375 -94 -1187 94
rect -1009 -94 -821 94
rect -643 -94 -455 94
rect -277 -94 -89 94
rect 89 -94 277 94
rect 455 -94 643 94
rect 821 -94 1009 94
rect 1187 -94 1375 94
rect 1553 -94 1741 94
<< locali >>
rect -1798 134 -1750 151
rect -1544 134 -1496 151
rect -1798 103 -1781 134
rect -1513 103 -1496 134
rect -1749 -94 -1741 94
rect -1553 -94 -1545 94
rect -1798 -134 -1781 -103
rect -1513 -134 -1496 -103
rect -1798 -151 -1750 -134
rect -1544 -151 -1496 -134
rect -1432 134 -1384 151
rect -1178 134 -1130 151
rect -1432 103 -1415 134
rect -1147 103 -1130 134
rect -1383 -94 -1375 94
rect -1187 -94 -1179 94
rect -1432 -134 -1415 -103
rect -1147 -134 -1130 -103
rect -1432 -151 -1384 -134
rect -1178 -151 -1130 -134
rect -1066 134 -1018 151
rect -812 134 -764 151
rect -1066 103 -1049 134
rect -781 103 -764 134
rect -1017 -94 -1009 94
rect -821 -94 -813 94
rect -1066 -134 -1049 -103
rect -781 -134 -764 -103
rect -1066 -151 -1018 -134
rect -812 -151 -764 -134
rect -700 134 -652 151
rect -446 134 -398 151
rect -700 103 -683 134
rect -415 103 -398 134
rect -651 -94 -643 94
rect -455 -94 -447 94
rect -700 -134 -683 -103
rect -415 -134 -398 -103
rect -700 -151 -652 -134
rect -446 -151 -398 -134
rect -334 134 -286 151
rect -80 134 -32 151
rect -334 103 -317 134
rect -49 103 -32 134
rect -285 -94 -277 94
rect -89 -94 -81 94
rect -334 -134 -317 -103
rect -49 -134 -32 -103
rect -334 -151 -286 -134
rect -80 -151 -32 -134
rect 32 134 80 151
rect 286 134 334 151
rect 32 103 49 134
rect 317 103 334 134
rect 81 -94 89 94
rect 277 -94 285 94
rect 32 -134 49 -103
rect 317 -134 334 -103
rect 32 -151 80 -134
rect 286 -151 334 -134
rect 398 134 446 151
rect 652 134 700 151
rect 398 103 415 134
rect 683 103 700 134
rect 447 -94 455 94
rect 643 -94 651 94
rect 398 -134 415 -103
rect 683 -134 700 -103
rect 398 -151 446 -134
rect 652 -151 700 -134
rect 764 134 812 151
rect 1018 134 1066 151
rect 764 103 781 134
rect 1049 103 1066 134
rect 813 -94 821 94
rect 1009 -94 1017 94
rect 764 -134 781 -103
rect 1049 -134 1066 -103
rect 764 -151 812 -134
rect 1018 -151 1066 -134
rect 1130 134 1178 151
rect 1384 134 1432 151
rect 1130 103 1147 134
rect 1415 103 1432 134
rect 1179 -94 1187 94
rect 1375 -94 1383 94
rect 1130 -134 1147 -103
rect 1415 -134 1432 -103
rect 1130 -151 1178 -134
rect 1384 -151 1432 -134
rect 1496 134 1544 151
rect 1750 134 1798 151
rect 1496 103 1513 134
rect 1781 103 1798 134
rect 1545 -94 1553 94
rect 1741 -94 1749 94
rect 1496 -134 1513 -103
rect 1781 -134 1798 -103
rect 1496 -151 1544 -134
rect 1750 -151 1798 -134
<< viali >>
rect -1741 -94 -1553 94
rect -1375 -94 -1187 94
rect -1009 -94 -821 94
rect -643 -94 -455 94
rect -277 -94 -89 94
rect 89 -94 277 94
rect 455 -94 643 94
rect 821 -94 1009 94
rect 1187 -94 1375 94
rect 1553 -94 1741 94
<< metal1 >>
rect -1747 94 -1547 97
rect -1747 -94 -1741 94
rect -1553 -94 -1547 94
rect -1747 -97 -1547 -94
rect -1381 94 -1181 97
rect -1381 -94 -1375 94
rect -1187 -94 -1181 94
rect -1381 -97 -1181 -94
rect -1015 94 -815 97
rect -1015 -94 -1009 94
rect -821 -94 -815 94
rect -1015 -97 -815 -94
rect -649 94 -449 97
rect -649 -94 -643 94
rect -455 -94 -449 94
rect -649 -97 -449 -94
rect -283 94 -83 97
rect -283 -94 -277 94
rect -89 -94 -83 94
rect -283 -97 -83 -94
rect 83 94 283 97
rect 83 -94 89 94
rect 277 -94 283 94
rect 83 -97 283 -94
rect 449 94 649 97
rect 449 -94 455 94
rect 643 -94 649 94
rect 449 -97 649 -94
rect 815 94 1015 97
rect 815 -94 821 94
rect 1009 -94 1015 94
rect 815 -97 1015 -94
rect 1181 94 1381 97
rect 1181 -94 1187 94
rect 1375 -94 1381 94
rect 1181 -97 1381 -94
rect 1547 94 1747 97
rect 1547 -94 1553 94
rect 1741 -94 1747 94
rect 1547 -97 1747 -94
<< properties >>
string FIXED_BBOX 1504 -142 1789 142
string gencell sky130_fd_pr__diode_pw2nd_05v5
string library sky130
string parameters w 2 l 2 area 4.0 peri 8.0 nx 10 ny 1 dummy 0 lmin 0.45 wmin 0.45 elc 1 erc 1 etc 1 ebc 1 doverlap 0 compatible {sky130_fd_pr__diode_pw2nd_05v5 sky130_fd_pr__diode_pw2nd_05v5_lvt  sky130_fd_pr__diode_pw2nd_05v5_nvt sky130_fd_pr__diode_pw2nd_11v0} full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
