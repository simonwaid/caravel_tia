magic
tech sky130A
magscale 1 2
timestamp 1647254192
<< pwell >>
rect -425 -1337 425 1337
<< nmos >>
rect -229 727 -29 1127
rect 29 727 229 1127
rect -229 109 -29 509
rect 29 109 229 509
rect -229 -509 -29 -109
rect 29 -509 229 -109
rect -229 -1127 -29 -727
rect 29 -1127 229 -727
<< ndiff >>
rect -287 1115 -229 1127
rect -287 739 -275 1115
rect -241 739 -229 1115
rect -287 727 -229 739
rect -29 1115 29 1127
rect -29 739 -17 1115
rect 17 739 29 1115
rect -29 727 29 739
rect 229 1115 287 1127
rect 229 739 241 1115
rect 275 739 287 1115
rect 229 727 287 739
rect -287 497 -229 509
rect -287 121 -275 497
rect -241 121 -229 497
rect -287 109 -229 121
rect -29 497 29 509
rect -29 121 -17 497
rect 17 121 29 497
rect -29 109 29 121
rect 229 497 287 509
rect 229 121 241 497
rect 275 121 287 497
rect 229 109 287 121
rect -287 -121 -229 -109
rect -287 -497 -275 -121
rect -241 -497 -229 -121
rect -287 -509 -229 -497
rect -29 -121 29 -109
rect -29 -497 -17 -121
rect 17 -497 29 -121
rect -29 -509 29 -497
rect 229 -121 287 -109
rect 229 -497 241 -121
rect 275 -497 287 -121
rect 229 -509 287 -497
rect -287 -739 -229 -727
rect -287 -1115 -275 -739
rect -241 -1115 -229 -739
rect -287 -1127 -229 -1115
rect -29 -739 29 -727
rect -29 -1115 -17 -739
rect 17 -1115 29 -739
rect -29 -1127 29 -1115
rect 229 -739 287 -727
rect 229 -1115 241 -739
rect 275 -1115 287 -739
rect 229 -1127 287 -1115
<< ndiffc >>
rect -275 739 -241 1115
rect -17 739 17 1115
rect 241 739 275 1115
rect -275 121 -241 497
rect -17 121 17 497
rect 241 121 275 497
rect -275 -497 -241 -121
rect -17 -497 17 -121
rect 241 -497 275 -121
rect -275 -1115 -241 -739
rect -17 -1115 17 -739
rect 241 -1115 275 -739
<< psubdiff >>
rect -389 1267 -293 1301
rect 293 1267 389 1301
rect -389 1205 -355 1267
rect 355 1205 389 1267
rect -389 -1267 -355 -1205
rect 355 -1267 389 -1205
rect -389 -1301 -293 -1267
rect 293 -1301 389 -1267
<< psubdiffcont >>
rect -293 1267 293 1301
rect -389 -1205 -355 1205
rect 355 -1205 389 1205
rect -293 -1301 293 -1267
<< poly >>
rect -229 1199 -29 1215
rect -229 1165 -213 1199
rect -45 1165 -29 1199
rect -229 1127 -29 1165
rect 29 1199 229 1215
rect 29 1165 45 1199
rect 213 1165 229 1199
rect 29 1127 229 1165
rect -229 689 -29 727
rect -229 655 -213 689
rect -45 655 -29 689
rect -229 639 -29 655
rect 29 689 229 727
rect 29 655 45 689
rect 213 655 229 689
rect 29 639 229 655
rect -229 581 -29 597
rect -229 547 -213 581
rect -45 547 -29 581
rect -229 509 -29 547
rect 29 581 229 597
rect 29 547 45 581
rect 213 547 229 581
rect 29 509 229 547
rect -229 71 -29 109
rect -229 37 -213 71
rect -45 37 -29 71
rect -229 21 -29 37
rect 29 71 229 109
rect 29 37 45 71
rect 213 37 229 71
rect 29 21 229 37
rect -229 -37 -29 -21
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect -229 -109 -29 -71
rect 29 -37 229 -21
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 29 -109 229 -71
rect -229 -547 -29 -509
rect -229 -581 -213 -547
rect -45 -581 -29 -547
rect -229 -597 -29 -581
rect 29 -547 229 -509
rect 29 -581 45 -547
rect 213 -581 229 -547
rect 29 -597 229 -581
rect -229 -655 -29 -639
rect -229 -689 -213 -655
rect -45 -689 -29 -655
rect -229 -727 -29 -689
rect 29 -655 229 -639
rect 29 -689 45 -655
rect 213 -689 229 -655
rect 29 -727 229 -689
rect -229 -1165 -29 -1127
rect -229 -1199 -213 -1165
rect -45 -1199 -29 -1165
rect -229 -1215 -29 -1199
rect 29 -1165 229 -1127
rect 29 -1199 45 -1165
rect 213 -1199 229 -1165
rect 29 -1215 229 -1199
<< polycont >>
rect -213 1165 -45 1199
rect 45 1165 213 1199
rect -213 655 -45 689
rect 45 655 213 689
rect -213 547 -45 581
rect 45 547 213 581
rect -213 37 -45 71
rect 45 37 213 71
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect -213 -581 -45 -547
rect 45 -581 213 -547
rect -213 -689 -45 -655
rect 45 -689 213 -655
rect -213 -1199 -45 -1165
rect 45 -1199 213 -1165
<< locali >>
rect -389 1267 -293 1301
rect 293 1267 389 1301
rect -389 1205 -355 1267
rect 355 1205 389 1267
rect -229 1165 -213 1199
rect -45 1165 -29 1199
rect 29 1165 45 1199
rect 213 1165 229 1199
rect -275 1115 -241 1131
rect -275 723 -241 739
rect -17 1115 17 1131
rect -17 723 17 739
rect 241 1115 275 1131
rect 241 723 275 739
rect -229 655 -213 689
rect -45 655 -29 689
rect 29 655 45 689
rect 213 655 229 689
rect -229 547 -213 581
rect -45 547 -29 581
rect 29 547 45 581
rect 213 547 229 581
rect -275 497 -241 513
rect -275 105 -241 121
rect -17 497 17 513
rect -17 105 17 121
rect 241 497 275 513
rect 241 105 275 121
rect -229 37 -213 71
rect -45 37 -29 71
rect 29 37 45 71
rect 213 37 229 71
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 213 -71 229 -37
rect -275 -121 -241 -105
rect -275 -513 -241 -497
rect -17 -121 17 -105
rect -17 -513 17 -497
rect 241 -121 275 -105
rect 241 -513 275 -497
rect -229 -581 -213 -547
rect -45 -581 -29 -547
rect 29 -581 45 -547
rect 213 -581 229 -547
rect -229 -689 -213 -655
rect -45 -689 -29 -655
rect 29 -689 45 -655
rect 213 -689 229 -655
rect -275 -739 -241 -723
rect -275 -1131 -241 -1115
rect -17 -739 17 -723
rect -17 -1131 17 -1115
rect 241 -739 275 -723
rect 241 -1131 275 -1115
rect -229 -1199 -213 -1165
rect -45 -1199 -29 -1165
rect 29 -1199 45 -1165
rect 213 -1199 229 -1165
rect -389 -1267 -355 -1205
rect 355 -1267 389 -1205
rect -389 -1301 -293 -1267
rect 293 -1301 389 -1267
<< viali >>
rect -213 1165 -45 1199
rect 45 1165 213 1199
rect -275 739 -241 1115
rect -17 739 17 1115
rect 241 739 275 1115
rect -213 655 -45 689
rect 45 655 213 689
rect -213 547 -45 581
rect 45 547 213 581
rect -275 121 -241 497
rect -17 121 17 497
rect 241 121 275 497
rect -213 37 -45 71
rect 45 37 213 71
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect -275 -497 -241 -121
rect -17 -497 17 -121
rect 241 -497 275 -121
rect -213 -581 -45 -547
rect 45 -581 213 -547
rect -213 -689 -45 -655
rect 45 -689 213 -655
rect -275 -1115 -241 -739
rect -17 -1115 17 -739
rect 241 -1115 275 -739
rect -213 -1199 -45 -1165
rect 45 -1199 213 -1165
<< metal1 >>
rect -225 1199 -33 1205
rect -225 1165 -213 1199
rect -45 1165 -33 1199
rect -225 1159 -33 1165
rect 33 1199 225 1205
rect 33 1165 45 1199
rect 213 1165 225 1199
rect 33 1159 225 1165
rect -281 1115 -235 1127
rect -281 739 -275 1115
rect -241 739 -235 1115
rect -281 727 -235 739
rect -23 1115 23 1127
rect -23 739 -17 1115
rect 17 739 23 1115
rect -23 727 23 739
rect 235 1115 281 1127
rect 235 739 241 1115
rect 275 739 281 1115
rect 235 727 281 739
rect -225 689 -33 695
rect -225 655 -213 689
rect -45 655 -33 689
rect -225 649 -33 655
rect 33 689 225 695
rect 33 655 45 689
rect 213 655 225 689
rect 33 649 225 655
rect -225 581 -33 587
rect -225 547 -213 581
rect -45 547 -33 581
rect -225 541 -33 547
rect 33 581 225 587
rect 33 547 45 581
rect 213 547 225 581
rect 33 541 225 547
rect -281 497 -235 509
rect -281 121 -275 497
rect -241 121 -235 497
rect -281 109 -235 121
rect -23 497 23 509
rect -23 121 -17 497
rect 17 121 23 497
rect -23 109 23 121
rect 235 497 281 509
rect 235 121 241 497
rect 275 121 281 497
rect 235 109 281 121
rect -225 71 -33 77
rect -225 37 -213 71
rect -45 37 -33 71
rect -225 31 -33 37
rect 33 71 225 77
rect 33 37 45 71
rect 213 37 225 71
rect 33 31 225 37
rect -225 -37 -33 -31
rect -225 -71 -213 -37
rect -45 -71 -33 -37
rect -225 -77 -33 -71
rect 33 -37 225 -31
rect 33 -71 45 -37
rect 213 -71 225 -37
rect 33 -77 225 -71
rect -281 -121 -235 -109
rect -281 -497 -275 -121
rect -241 -497 -235 -121
rect -281 -509 -235 -497
rect -23 -121 23 -109
rect -23 -497 -17 -121
rect 17 -497 23 -121
rect -23 -509 23 -497
rect 235 -121 281 -109
rect 235 -497 241 -121
rect 275 -497 281 -121
rect 235 -509 281 -497
rect -225 -547 -33 -541
rect -225 -581 -213 -547
rect -45 -581 -33 -547
rect -225 -587 -33 -581
rect 33 -547 225 -541
rect 33 -581 45 -547
rect 213 -581 225 -547
rect 33 -587 225 -581
rect -225 -655 -33 -649
rect -225 -689 -213 -655
rect -45 -689 -33 -655
rect -225 -695 -33 -689
rect 33 -655 225 -649
rect 33 -689 45 -655
rect 213 -689 225 -655
rect 33 -695 225 -689
rect -281 -739 -235 -727
rect -281 -1115 -275 -739
rect -241 -1115 -235 -739
rect -281 -1127 -235 -1115
rect -23 -739 23 -727
rect -23 -1115 -17 -739
rect 17 -1115 23 -739
rect -23 -1127 23 -1115
rect 235 -739 281 -727
rect 235 -1115 241 -739
rect 275 -1115 281 -739
rect 235 -1127 281 -1115
rect -225 -1165 -33 -1159
rect -225 -1199 -213 -1165
rect -45 -1199 -33 -1165
rect -225 -1205 -33 -1199
rect 33 -1165 225 -1159
rect 33 -1199 45 -1165
rect 213 -1199 225 -1165
rect 33 -1205 225 -1199
<< properties >>
string FIXED_BBOX -372 -1284 372 1284
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 1 m 4 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
