* SPICE3 file created from mpw5_submission_flat.ext - technology: sky130A

X0 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8 outd_0/InputRef tia_core_0/VM39D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X9 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X11 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X12 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X16 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X17 eigth_mirror_0/I_In isource_0/VM22D a_n35954_n3878# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X18 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X19 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X20 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X21 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X22 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X23 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X24 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X25 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X26 outd_0/outd_stage1_0/isource_out outd_0/InputRef outd_0/V_da1_N outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X27 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X28 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X29 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X30 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X31 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X32 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X33 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X34 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X35 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X36 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X37 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X38 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X39 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X40 cmirror_channel_0/VP outd_0/OutputP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X41 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X42 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X43 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X44 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X45 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X46 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X47 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X48 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X49 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X50 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X51 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X52 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X53 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X54 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X55 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X56 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X57 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X58 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X59 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X60 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X61 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X62 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X63 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X64 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X65 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X66 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X67 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X68 cmirror_channel_0/VP eigth_mirror_0/I_In a_n19500_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X69 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X70 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X71 cmirror_channel_0/VP outd_0/OutputP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X72 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X73 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X74 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X75 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X76 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X77 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X78 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X79 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X80 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X81 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X82 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X83 cmirror_channel_0/TIA_I_Bias1 a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X84 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X85 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X86 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X87 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X88 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X89 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X90 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X91 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X92 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X93 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X94 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X95 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X96 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X97 cmirror_channel_0/VN cmirror_channel_0/VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X98 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X99 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X100 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X101 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X102 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X103 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X104 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X105 isource_0/VM9D isource_0/VM9D isource_0/VM2D isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X106 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X107 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X108 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X109 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X110 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X111 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X112 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X113 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X114 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X115 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X116 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X117 a_n16800_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X118 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X119 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X120 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X121 cmirror_channel_0/VP eigth_mirror_0/I_In a_n22200_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X122 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X123 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X124 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X125 tia_core_0/VM39D cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM36D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X126 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X127 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X128 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X129 a_n5250_n3337# a_n5450_n3434# a_n5450_n3434# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X130 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X131 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X132 tia_core_0/VM31D outd_0/InputRef tia_core_0/VM39D tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X133 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X134 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X135 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X136 isource_0/VM2D isource_0/VM2D cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X137 cmirror_channel_0/VP isource_0/VM14D isource_0/VM12G isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X138 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X139 outd_0/InputRef tia_core_0/VM39D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X140 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X141 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X142 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X143 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X144 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X145 a_n35954_n3878# isource_0/VM22D eigth_mirror_0/I_In cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X146 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X147 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X148 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X149 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X150 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X151 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X152 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X153 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X154 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X155 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X156 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X157 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X158 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X159 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X160 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X161 a_n18150_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X162 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X163 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X164 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X165 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X166 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X167 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X168 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X169 tia_core_0/VM39D outd_0/InputRef tia_core_0/VM31D tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X170 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X171 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X172 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X173 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X174 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X175 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X176 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X177 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X178 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X179 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X180 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X181 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X182 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X183 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X184 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X185 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X186 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X187 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X188 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X189 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X190 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X191 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X192 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X193 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X194 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X195 isource_0/VM9D isource_0/VM9D isource_0/VM2D isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X196 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X197 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X198 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X199 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X200 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X201 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X202 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X203 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X204 tia_core_0/VM39D outd_0/InputRef tia_core_0/VM31D tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X205 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X206 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X207 cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM6D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X208 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X209 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X210 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X211 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X212 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X213 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X214 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X215 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X216 eigth_mirror_0/I_out_1 eigth_mirror_0/I_In a_n14100_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X217 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X218 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X219 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X220 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X221 a_n12750_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X222 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X223 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X224 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X225 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X226 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X227 eigth_mirror_0/I_out_5 eigth_mirror_0/I_In a_n19500_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X228 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X229 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X230 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X231 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X232 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X233 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X234 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X235 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X236 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X237 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X238 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X239 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X240 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X241 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X242 a_n19500_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X243 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X244 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X245 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X246 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X247 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X248 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X249 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X250 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X251 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X252 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X253 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X254 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X255 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X256 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X257 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X258 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X259 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X260 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X261 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X262 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X263 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X264 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X265 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X266 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X267 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X268 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X269 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X270 cmirror_channel_0/VP cmirror_channel_0/VN tia_core_0/VM31D cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X271 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X272 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X273 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X274 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X275 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X276 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X277 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X278 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X279 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X280 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X281 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X282 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X283 isource_0/VM3D isource_0/VM3G cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X284 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X285 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X286 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X287 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X288 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X289 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X290 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X291 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X292 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X293 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X294 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X295 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X296 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X297 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X298 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X299 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X300 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X301 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X302 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X303 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X304 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X305 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X306 isource_0/VM12G isource_0/VM14D cmirror_channel_0/VP isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X307 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X308 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X309 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X310 a_n25012_12290# isource_0/VM11D cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X311 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X312 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X313 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X314 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X315 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X316 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X317 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X318 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X319 cmirror_channel_0/VN cmirror_channel_0/I_in_channel a_n4672_n5100# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X320 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X321 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X322 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X323 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X324 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X325 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X326 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X327 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X328 outd_0/InputRef tia_core_0/VM39D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X329 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X330 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X331 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X332 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X333 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X334 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X335 a_n17034_6079# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X336 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X337 tia_core_0/Input outd_0/InputSignal tia_core_0/Out_2 tia_core_0/Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X338 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X339 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X340 a_n15450_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X341 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X342 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X343 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X344 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X345 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X346 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X347 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X348 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X349 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X350 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X351 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X352 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X353 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X354 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X355 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X356 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X357 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X358 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X359 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X360 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X361 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X362 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X363 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X364 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X365 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X366 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X367 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X368 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X369 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X370 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X371 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X372 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X373 outd_0/V_da2_N cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X374 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X375 tia_core_0/Input outd_0/InputSignal tia_core_0/Out_2 tia_core_0/Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X376 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X377 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X378 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X379 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X380 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X381 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X382 cmirror_channel_0/VN cmirror_channel_0/TIA_I_Bias1 sky130_fd_pr__cap_mim_m3_1 l=1.2e+07u w=1.5e+07u
X383 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X384 cmirror_channel_0/VP outd_0/OutputN cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X385 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X386 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X387 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X388 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X389 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X390 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X391 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X392 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X393 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X394 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X395 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X396 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X397 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X398 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X399 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X400 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X401 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X402 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X403 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X404 a_n17034_n701# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X405 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X406 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X407 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X408 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X409 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X410 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X411 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X412 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X413 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X414 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X415 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X416 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X417 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X418 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X419 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X420 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X421 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X422 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X423 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X424 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X425 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X426 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X427 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X428 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X429 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X430 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X431 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X432 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X433 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X434 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X435 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X436 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X437 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X438 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X439 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X440 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X441 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X442 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X443 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X444 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X445 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X446 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X447 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X448 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X449 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X450 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X451 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X452 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X453 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X454 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X455 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X456 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X457 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X458 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X459 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X460 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X461 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X462 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X463 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X464 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X465 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X466 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X467 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X468 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X469 tia_core_0/Input outd_0/InputSignal tia_core_0/Out_2 tia_core_0/Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X470 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X471 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X472 a_n5250_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X473 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X474 a_n20850_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X475 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X476 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X477 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X478 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X479 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X480 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X481 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X482 cmirror_channel_0/VP outd_0/V_da2_P cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X483 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X484 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X485 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X486 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X487 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X488 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X489 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X490 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X491 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X492 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X493 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X494 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X495 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X496 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X497 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X498 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X499 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X500 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X501 isource_0/VM9D isource_0/VM9D isource_0/VM2D isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X502 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X503 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X504 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X505 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X506 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X507 a_n11400_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X508 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X509 eigth_mirror_0/I_In isource_0/VM22D a_n35954_n3878# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X510 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X511 a_n19500_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X512 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X513 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X514 cmirror_channel_0/A_Out_I_Bias a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X515 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X516 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X517 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X518 tia_core_0/VM39D outd_0/InputRef tia_core_0/VM31D tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X519 isource_0/VM2D isource_0/VM9D isource_0/VM9D isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X520 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X521 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X522 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X523 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X524 cmirror_channel_0/VP outd_0/OutputN cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X525 cmirror_channel_0/VN cmirror_channel_0/VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X526 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X527 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X528 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X529 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X530 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X531 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X532 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X533 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X534 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X535 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X536 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X537 cmirror_channel_0/TIA_I_Bias1 a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X538 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X539 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X540 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X541 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X542 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X543 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X544 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X545 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X546 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X547 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X548 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X549 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X550 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X551 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X552 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X553 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X554 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X555 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X556 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X557 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X558 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X559 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X560 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X561 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X562 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X563 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X564 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X565 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X566 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X567 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X568 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X569 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X570 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X571 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X572 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X573 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X574 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X575 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X576 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X577 a_n17034_n701# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X578 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X579 cmirror_channel_0/VP isource_0/VM8D a_n17034_6079# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X580 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X581 cmirror_channel_0/VP eigth_mirror_0/I_In a_n20850_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X582 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X583 cmirror_channel_0/VN cmirror_channel_0/VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X584 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X585 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X586 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X587 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X588 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X589 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X590 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X591 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X592 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X593 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X594 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X595 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X596 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X597 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X598 cmirror_channel_0/VN isource_0/VM2D isource_0/VM2D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X599 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X600 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X601 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X602 cmirror_channel_0/VP outd_0/V_da2_P cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X603 outd_0/InputRef tia_core_0/VM39D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X604 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X605 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X606 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X607 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X608 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X609 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X610 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X611 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X612 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X613 cmirror_channel_0/VP eigth_mirror_0/I_In a_n22200_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X614 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X615 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X616 cmirror_channel_0/VP eigth_mirror_0/I_In a_n14100_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X617 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X618 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X619 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X620 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X621 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X622 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X623 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X624 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X625 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X626 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X627 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X628 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X629 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X630 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X631 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X632 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X633 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X634 cmirror_channel_0/VP outd_0/OutputP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X635 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X636 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X637 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X638 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X639 a_n35954_n3878# isource_0/VM22D eigth_mirror_0/I_In cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X640 outd_0/InputSignal tia_core_0/Input cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X641 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X642 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X643 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X644 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X645 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X646 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X647 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X648 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X649 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X650 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X651 outd_0/InputSignal tia_core_0/Input cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X652 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X653 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X654 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X655 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X656 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X657 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X658 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X659 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X660 a_n20850_n11957# eigth_mirror_0/I_In eigth_mirror_0/I_out_6 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X661 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X662 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X663 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X664 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X665 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X666 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X667 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X668 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X669 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X670 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X671 a_n5512_n5100# cmirror_channel_0/I_in_channel cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X672 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X673 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X674 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X675 a_n11400_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X676 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X677 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X678 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X679 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X680 cmirror_channel_0/TIA_I_Bias1 a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X681 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X682 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X683 a_n17034_n2971# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X684 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X685 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X686 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X687 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X688 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X689 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X690 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X691 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X692 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X693 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X694 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X695 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X696 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X697 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X698 a_n5450_n3434# cmirror_channel_0/I_in_channel a_n5512_n5100# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X699 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X700 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X701 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X702 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X703 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X704 tia_core_0/VM31D cmirror_channel_0/VN cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X705 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X706 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X707 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X708 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X709 tia_core_0/Out_2 outd_0/InputSignal tia_core_0/Input tia_core_0/Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X710 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X711 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X712 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X713 a_n12750_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X714 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X715 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X716 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X717 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X718 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X719 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X720 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X721 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X722 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X723 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X724 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X725 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X726 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X727 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X728 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X729 cmirror_channel_0/A_Out_I_Bias a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X730 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X731 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X732 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X733 cmirror_channel_0/VN isource_0/VM11D a_n25012_12290# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X734 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X735 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X736 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X737 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X738 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X739 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X740 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X741 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X742 outd_0/InputSignal tia_core_0/Input cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X743 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X744 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X745 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X746 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X747 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X748 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X749 outd_0/InputSignal tia_core_0/Input cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X750 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X751 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X752 tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__cap_var_lvt pd=0u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X753 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X754 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X755 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X756 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X757 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X758 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X759 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X760 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X761 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X762 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X763 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X764 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X765 cmirror_channel_0/VN isource_0/VM2D isource_0/VM2D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X766 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X767 eigth_mirror_0/I_out_1 eigth_mirror_0/I_In a_n14100_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X768 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X769 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X770 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X771 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X772 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X773 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X774 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X775 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X776 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X777 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X778 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X779 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X780 cmirror_channel_0/TIA_I_Bias1 a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X781 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X782 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X783 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X784 a_n14100_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X785 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X786 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X787 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X788 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X789 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X790 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X791 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X792 cmirror_channel_0/VN isource_0/VM2D isource_0/VM2D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X793 tia_core_0/VM31D outd_0/InputRef tia_core_0/VM39D tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X794 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X795 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X796 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X797 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X798 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X799 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X800 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X801 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X802 cmirror_channel_0/VN cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM36D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X803 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X804 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X805 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X806 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X807 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X808 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X809 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X810 outd_0/V_da1_N outd_0/InputRef outd_0/outd_stage1_0/isource_out outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X811 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X812 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X813 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X814 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X815 a_n15450_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X816 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X817 a_17268_7820# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X818 outd_0/V_da2_N cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X819 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X820 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X821 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X822 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X823 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X824 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X825 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X826 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X827 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X828 cmirror_channel_0/A_Out_I_Bias a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X829 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X830 cmirror_channel_0/VN isource_0/VM11D a_n25012_12290# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X831 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X832 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X833 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X834 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X835 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X836 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X837 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X838 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X839 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X840 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X841 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X842 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X843 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X844 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X845 outd_0/InputSignal tia_core_0/Input cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X846 isource_0/VM12G isource_0/VM14D cmirror_channel_0/VP isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X847 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X848 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X849 cmirror_channel_0/VP eigth_mirror_0/I_In a_n19500_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X850 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X851 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X852 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X853 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X854 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X855 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X856 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X857 cmirror_channel_0/VP isource_0/VM8D a_n17034_n2971# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X858 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X859 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X860 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X861 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X862 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X863 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X864 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X865 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X866 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X867 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X868 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X869 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X870 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X871 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X872 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X873 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X874 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X875 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X876 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X877 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X878 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X879 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X880 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X881 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X882 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X883 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X884 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X885 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X886 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X887 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X888 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X889 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X890 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X891 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X892 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X893 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X894 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X895 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X896 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X897 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X898 cmirror_channel_0/VP eigth_mirror_0/I_In a_n16800_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X899 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X900 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X901 cmirror_channel_0/A_Out_I_Bias a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X902 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X903 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X904 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X905 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X906 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X907 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X908 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X909 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X910 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X911 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X912 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X913 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X914 cmirror_channel_0/VP eigth_mirror_0/I_In a_n22200_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X915 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X916 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X917 cmirror_channel_0/TIA_I_Bias1 a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X918 isource_0/VM8D isource_0/VM9D isource_0/VM11D isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X919 cmirror_channel_0/VP outd_0/OutputN cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X920 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X921 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X922 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X923 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X924 cmirror_channel_0/VP eigth_mirror_0/I_In a_n15450_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X925 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X926 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X927 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X928 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X929 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X930 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X931 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X932 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X933 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X934 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X935 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X936 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X937 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X938 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X939 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X940 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X941 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X942 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X943 cmirror_channel_0/VP a_n5450_n3434# a_n5250_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X944 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X945 cmirror_channel_0/VP eigth_mirror_0/I_In a_n20850_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X946 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X947 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X948 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X949 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X950 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X951 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X952 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X953 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X954 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X955 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X956 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X957 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X958 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X959 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X960 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X961 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X962 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X963 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X964 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X965 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X966 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X967 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X968 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X969 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X970 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X971 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X972 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X973 cmirror_channel_0/VN isource_0/VM2D isource_0/VM2D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X974 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X975 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X976 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X977 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X978 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X979 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X980 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X981 a_n19500_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X982 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X983 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X984 cmirror_channel_0/VP isource_0/VM8D a_n17034_n2971# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X985 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X986 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X987 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X988 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X989 isource_0/VM3D a_n35954_n3878# isource_0/VM22D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X990 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X991 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X992 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X993 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X994 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X995 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X996 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X997 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X998 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X999 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1000 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1001 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1002 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1003 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1004 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1005 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1006 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1007 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1008 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1009 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1010 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1011 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1012 a_n15450_n11957# eigth_mirror_0/I_In eigth_mirror_0/I_out_2 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1013 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1014 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1015 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1016 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1017 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1018 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1019 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1020 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1021 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1022 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1023 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1024 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1025 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1026 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1027 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1028 cmirror_channel_0/A_Out_I_Bias a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1029 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1030 isource_0/VM8D isource_0/VM9D isource_0/VM11D isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1031 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1032 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1033 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1034 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1035 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1036 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1037 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1038 cmirror_channel_0/VP eigth_mirror_0/I_In a_n11400_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1039 cmirror_channel_0/TIA_I_Bias1 a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1040 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1041 cmirror_channel_0/VN cmirror_channel_0/I_in_channel a_n4672_n5100# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1042 cmirror_channel_0/VP outd_0/OutputN cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1043 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1044 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1045 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1046 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1047 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1048 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1049 cmirror_channel_0/VP outd_0/OutputP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1050 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1051 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1052 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1053 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1054 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1055 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1056 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1057 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1058 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1059 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1060 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1061 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1062 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1063 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1064 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1065 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1066 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1067 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1068 eigth_mirror_0/I_In isource_0/VM22D a_n35954_n3878# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1069 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1070 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1071 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1072 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1073 cmirror_channel_0/VN cmirror_channel_0/VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1074 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1075 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1076 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1077 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1078 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1079 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1080 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1081 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1082 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1083 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1084 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1085 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1086 isource_0/VM3D a_n35954_n3878# isource_0/VM22D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1087 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1088 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1089 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1090 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1091 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1092 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1093 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1094 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1095 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1096 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1097 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1098 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1099 tia_core_0/Input outd_0/InputSignal tia_core_0/Out_2 tia_core_0/Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1100 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1101 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1102 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1103 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1104 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1105 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1106 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1107 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1108 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1109 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1110 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1111 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1112 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1113 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1114 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1115 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1116 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1117 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1118 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1119 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1120 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1121 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1122 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1123 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1124 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1125 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1126 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1127 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1128 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1129 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1130 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1131 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1132 a_n17034_n701# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1133 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1134 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1135 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1136 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1137 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1138 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1139 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1140 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1141 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1142 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1143 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1144 a_n15450_n11957# eigth_mirror_0/I_In eigth_mirror_0/I_out_2 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1145 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1146 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1147 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1148 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1149 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1150 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1151 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1152 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1153 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1154 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1155 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1156 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1157 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1158 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1159 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1160 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1161 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1162 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1163 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1164 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1165 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1166 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1167 a_n18994_26# a_n19524_2458# cmirror_channel_0/VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X1168 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1169 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1170 a_n14100_n11957# eigth_mirror_0/I_In eigth_mirror_0/I_out_1 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1171 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1172 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1173 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1174 cmirror_channel_0/VP outd_0/OutputP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1175 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1176 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1177 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1178 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1179 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1180 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1181 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1182 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1183 tia_core_0/VM39D cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM36D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1184 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1185 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1186 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1187 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1188 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1189 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1190 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1191 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1192 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1193 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1194 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1195 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1196 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1197 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1198 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1199 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1200 isource_0/VM11D isource_0/VM9D isource_0/VM8D isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1201 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1202 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1203 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1204 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1205 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1206 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1207 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1208 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1209 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1210 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1211 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1212 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1213 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1214 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1215 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1216 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1217 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1218 outd_0/V_da1_P outd_0/InputSignal outd_0/outd_stage1_0/isource_out outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1219 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1220 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1221 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1222 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1223 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1224 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1225 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1226 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1227 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1228 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1229 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1230 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1231 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1232 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1233 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1234 cmirror_channel_0/VN cmirror_channel_0/TIA_I_Bias1 sky130_fd_pr__cap_mim_m3_1 l=1.2e+07u w=1.5e+07u
X1235 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1236 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1237 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1238 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1239 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1240 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1241 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1242 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1243 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1244 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1245 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1246 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1247 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1248 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1249 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1250 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1251 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1252 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1253 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1254 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1255 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1256 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1257 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1258 cmirror_channel_0/VN cmirror_channel_0/VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1259 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1260 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1261 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1262 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1263 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1264 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1265 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1266 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1267 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1268 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1269 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1270 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1271 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1272 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1273 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1274 cmirror_channel_0/TIA_I_Bias1 a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1275 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1276 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1277 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1278 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1279 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1280 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1281 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1282 outd_0/InputRef tia_core_0/VM39D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1283 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1284 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1285 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1286 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1287 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1288 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1289 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1290 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1291 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1292 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1293 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1294 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1295 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1296 outd_0/OutputN cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1297 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1298 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1299 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1300 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1301 cmirror_channel_0/VP eigth_mirror_0/I_In a_n16800_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1302 isource_0/VM22D a_n35954_n3878# isource_0/VM3D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1303 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1304 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1305 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1306 a_n35954_n3878# isource_0/VM22D eigth_mirror_0/I_In cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1307 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1308 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1309 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1310 outd_0/InputRef tia_core_0/VM39D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1311 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1312 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1313 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1314 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1315 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1316 cmirror_channel_0/VP eigth_mirror_0/I_In a_n18150_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1317 tia_core_0/Input cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM5D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1318 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1319 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1320 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1321 a_n17034_n701# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1322 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1323 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1324 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1325 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1326 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1327 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1328 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1329 a_n22200_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1330 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1331 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1332 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1333 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1334 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1335 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1336 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1337 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1338 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1339 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1340 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1341 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1342 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1343 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1344 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1345 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1346 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1347 cmirror_channel_0/VP cmirror_channel_0/VN tia_core_0/Out_2 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1348 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1349 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1350 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1351 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1352 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1353 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1354 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1355 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1356 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1357 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1358 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1359 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1360 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1361 cmirror_channel_0/VN cmirror_channel_0/VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1362 outd_0/InputSignal tia_core_0/Input cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1363 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1364 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1365 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1366 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1367 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1368 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1369 isource_0/VM11D isource_0/VM9D isource_0/VM8D isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1370 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1371 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1372 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1373 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1374 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1375 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1376 isource_0/VM22D a_n35954_n3878# isource_0/VM3D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1377 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1378 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1379 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1380 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1381 cmirror_channel_0/VP isource_0/VM8D a_n17034_8339# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1382 a_n16464_n6284# a_n15934_n3852# cmirror_channel_0/VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X1383 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1384 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1385 outd_0/V_da1_P outd_0/InputSignal outd_0/outd_stage1_0/isource_out outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1386 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1387 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1388 a_n17034_6079# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1389 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1390 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1391 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1392 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1393 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1394 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1395 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1396 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1397 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1398 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1399 cmirror_channel_0/VP eigth_mirror_0/I_In a_n22200_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1400 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1401 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1402 cmirror_channel_0/VP eigth_mirror_0/I_In a_n14100_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1403 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1404 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1405 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1406 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1407 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1408 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1409 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1410 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1411 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1412 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1413 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1414 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1415 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1416 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1417 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1418 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1419 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1420 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1421 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1422 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1423 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1424 cmirror_channel_0/VP eigth_mirror_0/I_In a_n20850_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1425 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1426 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1427 cmirror_channel_0/VP eigth_mirror_0/I_In a_n12750_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1428 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1429 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1430 tia_core_0/VM6D cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1431 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1432 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1433 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1434 outd_0/outd_stage1_0/isource_out outd_0/InputSignal outd_0/V_da1_P outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1435 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1436 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1437 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1438 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1439 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1440 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1441 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1442 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1443 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1444 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1445 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1446 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1447 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1448 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1449 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1450 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1451 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1452 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1453 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1454 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1455 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1456 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1457 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1458 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1459 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1460 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1461 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1462 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1463 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1464 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1465 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1466 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1467 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1468 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1469 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1470 isource_0/VM22D a_n35954_n3878# isource_0/VM3D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1471 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1472 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1473 cmirror_channel_0/A_Out_I_Bias a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1474 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1475 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1476 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1477 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1478 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1479 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1480 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1481 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1482 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1483 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1484 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1485 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1486 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1487 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1488 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1489 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1490 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1491 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1492 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1493 isource_0/VM9D isource_0/VM9D isource_0/VM2D isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1494 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1495 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1496 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1497 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1498 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1499 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1500 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1501 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1502 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1503 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1504 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1505 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1506 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1507 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1508 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1509 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1510 a_n17034_n701# isource_0/VM8D isource_0/VM14D cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X1511 a_n17034_n701# isource_0/VM8D isource_0/VM14D cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X1512 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1513 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1514 cmirror_channel_0/VP eigth_mirror_0/I_In a_n11400_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1515 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1516 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1517 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1518 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1519 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1520 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1521 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1522 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1523 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1524 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1525 outd_0/InputRef tia_core_0/VM39D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1526 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1527 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1528 outd_0/InputRef tia_core_0/VM39D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1529 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1530 a_n21114_26# a_n21644_2458# cmirror_channel_0/VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X1531 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1532 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1533 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1534 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1535 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1536 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1537 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1538 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1539 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1540 outd_0/V_da1_N outd_0/InputRef outd_0/outd_stage1_0/isource_out outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1541 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1542 a_n17034_8339# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1543 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1544 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1545 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1546 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1547 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1548 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1549 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1550 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1551 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1552 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1553 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1554 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1555 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1556 tia_core_0/VM5D cmirror_channel_0/TIA_I_Bias1 tia_core_0/Input cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1557 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1558 isource_0/VM22D a_n35954_n3878# isource_0/VM3D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1559 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1560 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1561 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1562 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1563 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1564 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1565 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1566 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1567 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1568 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1569 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1570 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1571 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1572 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1573 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1574 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1575 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1576 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1577 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1578 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1579 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1580 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1581 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1582 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1583 cmirror_channel_0/VP outd_0/OutputP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1584 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1585 cmirror_channel_0/A_Out_I_Bias a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1586 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1587 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1588 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1589 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1590 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1591 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1592 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1593 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1594 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1595 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1596 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1597 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1598 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1599 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1600 tia_core_0/VM39D outd_0/InputRef tia_core_0/VM31D tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1601 cmirror_channel_0/VP outd_0/V_da2_N cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1602 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1603 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1604 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1605 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1606 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1607 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1608 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1609 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1610 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1611 tia_core_0/VM39D cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM36D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1612 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1613 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1614 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1615 cmirror_channel_0/VP isource_0/VM8D a_n17034_6079# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1616 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1617 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1618 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1619 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1620 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1621 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1622 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1623 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1624 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1625 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1626 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1627 isource_0/VM12G isource_0/VM14D cmirror_channel_0/VP isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1628 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1629 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1630 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1631 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1632 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1633 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1634 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1635 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1636 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1637 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1638 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1639 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1640 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1641 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1642 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1643 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1644 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1645 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1646 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1647 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1648 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1649 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1650 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1651 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1652 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1653 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1654 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1655 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1656 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1657 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1658 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1659 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1660 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1661 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1662 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1663 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1664 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1665 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1666 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1667 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1668 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1669 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1670 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1671 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1672 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1673 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1674 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1675 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1676 isource_0/VM11D isource_0/VM9D isource_0/VM8D isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1677 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1678 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1679 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1680 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1681 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1682 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1683 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1684 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1685 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1686 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1687 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1688 a_n17034_n701# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1689 a_n18150_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1690 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1691 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1692 a_n17034_n701# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1693 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1694 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1695 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1696 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1697 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1698 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1699 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1700 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1701 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1702 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1703 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1704 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1705 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1706 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1707 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1708 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1709 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1710 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1711 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1712 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1713 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1714 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1715 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1716 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1717 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1718 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1719 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1720 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1721 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1722 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1723 a_n17034_n701# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1724 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1725 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1726 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1727 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1728 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1729 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1730 cmirror_channel_0/VP outd_0/OutputP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1731 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1732 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1733 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1734 tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__cap_var_lvt pd=0u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X1735 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1736 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1737 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1738 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1739 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1740 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1741 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1742 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1743 tia_core_0/Out_2 cmirror_channel_0/VN cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1744 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1745 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1746 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1747 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1748 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1749 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1750 outd_0/InputRef tia_core_0/VM39D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1751 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1752 cmirror_channel_0/VP eigth_mirror_0/I_In a_n15450_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1753 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1754 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1755 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1756 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1757 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1758 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1759 eigth_mirror_0/I_out_7 eigth_mirror_0/I_In a_n22200_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1760 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1761 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1762 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1763 a_n20850_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1764 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1765 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1766 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1767 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1768 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1769 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1770 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1771 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1772 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1773 cmirror_channel_0/VN cmirror_channel_0/I_in_channel a_n5512_n5100# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1774 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1775 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1776 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1777 cmirror_channel_0/VN cmirror_channel_0/I_in_channel a_n4672_n5100# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1778 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1779 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1780 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1781 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1782 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1783 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1784 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1785 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1786 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1787 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1788 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1789 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1790 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1791 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1792 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1793 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1794 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1795 cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM6D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1796 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1797 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1798 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1799 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1800 cmirror_channel_0/VP eigth_mirror_0/I_In a_n16800_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1801 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1802 isource_0/VM3D a_n35954_n3878# isource_0/VM22D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1803 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1804 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1805 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1806 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1807 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1808 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1809 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1810 tia_core_0/VM36D cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM39D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1811 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1812 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1813 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1814 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1815 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1816 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1817 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1818 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1819 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1820 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1821 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1822 cmirror_channel_0/VN tia_core_0/Disable_TIA cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1823 cmirror_channel_0/VP eigth_mirror_0/I_In a_n18150_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1824 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1825 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1826 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1827 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1828 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1829 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1830 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1831 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1832 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1833 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1834 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1835 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1836 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1837 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1838 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1839 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1840 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1841 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1842 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1843 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1844 isource_0/VM8D isource_0/VM9D isource_0/VM11D isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1845 tia_core_0/VM39D outd_0/InputRef tia_core_0/VM31D tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1846 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1847 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1848 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1849 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1850 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1851 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1852 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1853 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1854 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1855 a_n16800_n11957# eigth_mirror_0/I_In eigth_mirror_0/I_out_3 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1856 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1857 cmirror_channel_0/VP eigth_mirror_0/I_In a_n11400_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1858 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1859 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1860 outd_0/outd_stage1_0/isource_out outd_0/InputRef outd_0/V_da1_N outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1861 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1862 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1863 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1864 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1865 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1866 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1867 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1868 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1869 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1870 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1871 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1872 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1873 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1874 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1875 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1876 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1877 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1878 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1879 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1880 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1881 a_n35954_n3878# isource_0/VM22D eigth_mirror_0/I_In cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1882 cmirror_channel_0/VP eigth_mirror_0/I_In a_n12750_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1883 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1884 isource_0/VM3D a_n35954_n3878# isource_0/VM22D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1885 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1886 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1887 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1888 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1889 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1890 outd_0/InputRef tia_core_0/VM39D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1891 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1892 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1893 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1894 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1895 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1896 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1897 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1898 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1899 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1900 outd_0/InputSignal tia_core_0/Input cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1901 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1902 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1903 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1904 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1905 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1906 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1907 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1908 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1909 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1910 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1911 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1912 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1913 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1914 tia_core_0/VM39D outd_0/InputRef tia_core_0/VM31D tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1915 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1916 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1917 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X1918 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1919 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1920 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1921 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1922 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1923 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1924 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1925 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1926 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1927 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1928 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1929 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1930 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1931 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1932 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1933 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1934 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1935 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1936 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1937 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1938 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1939 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1940 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1941 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1942 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1943 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1944 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1945 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1946 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1947 tia_core_0/VM5D cmirror_channel_0/TIA_I_Bias1 tia_core_0/Input cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1948 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1949 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1950 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1951 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1952 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1953 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1954 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1955 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1956 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1957 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1958 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1959 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1960 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1961 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1962 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1963 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1964 tia_core_0/VM31D cmirror_channel_0/VN cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1965 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1966 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1967 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1968 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1969 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1970 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1971 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1972 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1973 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1974 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1975 tia_core_0/VM31D outd_0/InputRef tia_core_0/VM39D tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1976 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1977 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1978 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1979 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1980 tia_core_0/Out_2 outd_0/InputSignal tia_core_0/Input tia_core_0/Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1981 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1982 cmirror_channel_0/VP cmirror_channel_0/VN tia_core_0/VM31D cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1983 cmirror_channel_0/VP isource_0/VM14D isource_0/VM12G isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1984 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1985 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1986 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1987 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1988 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1989 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1990 a_n20850_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1991 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1992 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1993 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X1994 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1995 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1996 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1997 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1998 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1999 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2000 outd_0/InputSignal tia_core_0/Input cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2001 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2002 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2003 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2004 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2005 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2006 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2007 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2008 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2009 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2010 outd_0/outd_stage1_0/isource_out outd_0/InputSignal outd_0/V_da1_P outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2011 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2012 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2013 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2014 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2015 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2016 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2017 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2018 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2019 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2020 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2021 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2022 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2023 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2024 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2025 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2026 isource_0/VM2D isource_0/VM2D cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X2027 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2028 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X2029 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2030 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2031 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2032 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2033 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2034 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2035 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2036 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2037 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2038 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2039 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2040 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2041 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2042 outd_0/OutputN cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2043 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2044 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2045 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2046 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2047 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2048 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2049 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2050 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2051 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X2052 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2053 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2054 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2055 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2056 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2057 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2058 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2059 cmirror_channel_0/VP outd_0/OutputN cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2060 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2061 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2062 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2063 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2064 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2065 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2066 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2067 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2068 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2069 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2070 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2071 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2072 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2073 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2074 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2075 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2076 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2077 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2078 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2079 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2080 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2081 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2082 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2083 a_n6352_n5100# cmirror_channel_0/I_in_channel cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2084 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2085 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2086 outd_0/V_da1_N outd_0/InputRef outd_0/outd_stage1_0/isource_out outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2087 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2088 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2089 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2090 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2091 eigth_mirror_0/I_out_4 eigth_mirror_0/I_In a_n18150_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2092 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2093 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2094 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2095 tia_core_0/Out_2 outd_0/InputSignal tia_core_0/Input tia_core_0/Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2096 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2097 a_n17034_8339# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2098 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2099 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2100 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2101 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2102 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2103 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2104 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2105 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2106 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2107 eigth_mirror_0/I_In isource_0/VM22D a_n35954_n3878# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2108 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2109 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2110 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2111 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2112 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2113 cmirror_channel_0/I_in_channel cmirror_channel_0/I_in_channel a_n6352_n5100# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2114 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2115 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2116 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2117 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2118 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2119 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2120 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2121 isource_0/VM11D isource_0/VM9D isource_0/VM8D isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2122 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2123 a_n5250_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2124 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2125 cmirror_channel_0/VP eigth_mirror_0/I_In a_n18150_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2126 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2127 tia_core_0/VM5D cmirror_channel_0/TIA_I_Bias1 tia_core_0/Input cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2128 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2129 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2130 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2131 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2132 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2133 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2134 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2135 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2136 cmirror_channel_0/VP eigth_mirror_0/I_In a_n22200_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2137 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2138 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2139 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2140 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2141 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2142 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2143 cmirror_channel_0/VP outd_0/OutputP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2144 cmirror_channel_0/VN cmirror_channel_0/VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2145 a_n17034_n701# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2146 a_n5250_n3337# a_n5450_n3434# a_n5450_n3434# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2147 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2148 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2149 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2150 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2151 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2152 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2153 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2154 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2155 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2156 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2157 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2158 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2159 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2160 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2161 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2162 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2163 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2164 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2165 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2166 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2167 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2168 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2169 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2170 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2171 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2172 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2173 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2174 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2175 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2176 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2177 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2178 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2179 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2180 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2181 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2182 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2183 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2184 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2185 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2186 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2187 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2188 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2189 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2190 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2191 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2192 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2193 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2194 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2195 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2196 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2197 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2198 outd_0/V_da1_N outd_0/InputRef outd_0/outd_stage1_0/isource_out outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2199 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2200 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2201 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2202 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2203 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2204 outd_0/outd_stage1_0/isource_out outd_0/InputSignal outd_0/V_da1_P outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2205 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2206 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2207 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2208 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2209 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2210 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2211 tia_core_0/VM31D outd_0/InputRef tia_core_0/VM39D tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2212 tia_core_0/Out_2 outd_0/InputSignal tia_core_0/Input tia_core_0/Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2213 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2214 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2215 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X2216 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2217 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2218 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2219 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2220 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2221 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2222 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2223 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2224 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2225 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2226 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2227 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2228 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2229 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2230 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2231 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2232 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2233 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2234 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2235 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2236 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2237 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2238 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2239 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2240 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2241 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2242 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2243 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2244 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2245 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2246 a_n20850_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2247 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2248 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2249 a_n12750_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2250 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2251 a_n17034_n701# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2252 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2253 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2254 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2255 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2256 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2257 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2258 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2259 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2260 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X2261 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2262 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2263 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2264 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2265 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2266 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2267 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2268 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2269 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2270 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2271 outd_0/OutputN cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2272 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2273 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2274 a_n17034_n701# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2275 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2276 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2277 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2278 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2279 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2280 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2281 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2282 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2283 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2284 isource_0/VM2D isource_0/VM2D cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X2285 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2286 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2287 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X2288 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2289 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2290 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2291 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2292 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2293 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2294 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2295 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2296 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2297 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2298 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2299 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2300 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2301 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2302 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2303 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2304 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2305 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2306 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2307 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2308 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2309 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2310 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2311 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2312 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2313 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2314 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2315 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2316 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2317 eigth_mirror_0/I_out_7 eigth_mirror_0/I_In a_n22200_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2318 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2319 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2320 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2321 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2322 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2323 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2324 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2325 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2326 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2327 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2328 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2329 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2330 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2331 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2332 tia_core_0/Input outd_0/InputSignal tia_core_0/Out_2 tia_core_0/Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2333 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2334 cmirror_channel_0/VP isource_0/VM8D a_n17034_8339# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2335 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2336 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2337 outd_0/V_da1_P outd_0/InputSignal outd_0/outd_stage1_0/isource_out outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2338 cmirror_channel_0/VP a_n5450_n3434# a_n5250_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2339 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2340 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2341 a_n22200_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2342 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2343 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2344 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2345 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2346 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2347 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2348 cmirror_channel_0/VP eigth_mirror_0/I_In a_n11400_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2349 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2350 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2351 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2352 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2353 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2354 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2355 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2356 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2357 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2358 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2359 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2360 a_n25012_12290# isource_0/VM11D cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X2361 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2362 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2363 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2364 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2365 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2366 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2367 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2368 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2369 outd_0/V_da2_P cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2370 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2371 outd_0/OutputN cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2372 outd_0/outd_stage1_0/isource_out outd_0/InputRef outd_0/V_da1_N outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2373 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2374 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2375 cmirror_channel_0/VP tia_core_0/VM28D sky130_fd_pr__cap_mim_m3_2 l=1.8e+07u w=2.5e+07u
X2376 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2377 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2378 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2379 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2380 cmirror_channel_0/VP eigth_mirror_0/I_In a_n12750_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2381 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2382 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2383 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2384 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2385 cmirror_channel_0/VP isource_0/VM11D a_n25012_12290# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X2386 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2387 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2388 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2389 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2390 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2391 a_n15450_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2392 tia_core_0/Input cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM5D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2393 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2394 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2395 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2396 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2397 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2398 a_n5250_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2399 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2400 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2401 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2402 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2403 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2404 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2405 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2406 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2407 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2408 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2409 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2410 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2411 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2412 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2413 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2414 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2415 cmirror_channel_0/VN isource_0/VM3G isource_0/VM3D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X2416 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2417 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2418 cmirror_channel_0/VP tia_core_0/Disable_TIA tia_core_0/Disable_TIA_B cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=1e+06u
X2419 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2420 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2421 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2422 outd_0/V_da1_N cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
X2423 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2424 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2425 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2426 outd_0/OutputP cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2427 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2428 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2429 cmirror_channel_0/VN cmirror_channel_0/I_in_channel a_n6352_n5100# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2430 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2431 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2432 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2433 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2434 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2435 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2436 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2437 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2438 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2439 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2440 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2441 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2442 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2443 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2444 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2445 tia_core_0/VM39D cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM36D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2446 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2447 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2448 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2449 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2450 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2451 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2452 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2453 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2454 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2455 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X2456 cmirror_channel_0/VP isource_0/VM14D isource_0/VM12G isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2457 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2458 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2459 tia_core_0/Input outd_0/InputSignal tia_core_0/Out_2 tia_core_0/Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2460 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2461 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2462 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2463 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2464 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2465 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2466 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2467 isource_0/VM9D isource_0/VM9D isource_0/VM2D isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2468 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2469 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2470 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2471 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2472 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2473 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2474 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2475 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2476 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2477 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2478 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2479 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2480 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2481 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2482 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2483 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2484 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2485 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2486 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2487 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2488 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2489 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2490 a_n25012_12290# isource_0/VM11D cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X2491 outd_0/InputRef tia_core_0/VM39D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2492 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2493 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2494 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2495 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2496 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2497 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2498 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2499 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2500 a_n17034_n2971# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2501 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2502 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2503 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2504 cmirror_channel_0/VN cmirror_channel_0/I_in_channel a_n5512_n5100# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2505 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2506 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2507 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2508 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2509 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2510 tia_core_0/Input outd_0/InputSignal tia_core_0/Out_2 tia_core_0/Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2511 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2512 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2513 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2514 outd_0/V_da2_P cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2515 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2516 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2517 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2518 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2519 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2520 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2521 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2522 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2523 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2524 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2525 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2526 isource_0/VM11D isource_0/VM9D isource_0/VM8D isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2527 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2528 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2529 cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM6D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2530 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2531 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2532 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2533 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2534 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2535 outd_0/OutputP cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2536 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2537 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2538 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2539 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2540 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2541 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2542 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2543 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2544 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2545 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2546 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2547 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2548 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2549 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2550 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2551 a_n19500_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2552 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2553 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2554 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2555 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2556 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2557 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2558 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2559 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2560 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2561 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2562 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2563 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2564 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2565 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2566 cmirror_channel_0/VP isource_0/VM14D isource_0/VM12G isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2567 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2568 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2569 tia_core_0/VM6D cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2570 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2571 a_n15450_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2572 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2573 cmirror_channel_0/VP a_n5450_n3434# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2574 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2575 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2576 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2577 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2578 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2579 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2580 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2581 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2582 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2583 tia_core_0/VM31D outd_0/InputRef tia_core_0/VM39D tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2584 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2585 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2586 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2587 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2588 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2589 outd_0/outd_stage1_0/isource_out outd_0/InputSignal outd_0/V_da1_P outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2590 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2591 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2592 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2593 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2594 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2595 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2596 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2597 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2598 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2599 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2600 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2601 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2602 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2603 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2604 a_n14100_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2605 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2606 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2607 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2608 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2609 tia_core_0/Out_2 cmirror_channel_0/VN cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2610 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2611 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2612 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2613 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X2614 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2615 outd_0/outd_stage1_0/isource_out outd_0/InputSignal outd_0/V_da1_P outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2616 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2617 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2618 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2619 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2620 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2621 a_n4672_n5100# cmirror_channel_0/I_in_channel cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2622 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2623 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2624 tia_core_0/Input outd_0/InputSignal tia_core_0/Out_2 tia_core_0/Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2625 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2626 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2627 tia_core_0/VM6D cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2628 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2629 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2630 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2631 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2632 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2633 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2634 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2635 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2636 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2637 a_n17034_6079# isource_0/VM8D isource_0/VM8D cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X2638 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2639 isource_0/VM12G isource_0/VM14D cmirror_channel_0/VP isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2640 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2641 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2642 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2643 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X2644 cmirror_channel_0/VP eigth_mirror_0/I_In a_n18150_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2645 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2646 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2647 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2648 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2649 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2650 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2651 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2652 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2653 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2654 cmirror_channel_0/VP outd_0/OutputN cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2655 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2656 tia_core_0/VM39D outd_0/InputRef tia_core_0/VM31D tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2657 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2658 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2659 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2660 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2661 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2662 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2663 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2664 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2665 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2666 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2667 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2668 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2669 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2670 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2671 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2672 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2673 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2674 outd_0/OutputP cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2675 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2676 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2677 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2678 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2679 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2680 cmirror_channel_0/I_in_channel eigth_mirror_0/I_In a_n12750_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2681 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2682 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2683 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2684 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2685 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2686 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2687 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2688 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2689 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2690 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2691 eigth_mirror_0/I_out_4 eigth_mirror_0/I_In a_n18150_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2692 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2693 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2694 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2695 outd_0/V_da1_N outd_0/InputRef outd_0/outd_stage1_0/isource_out outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2696 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2697 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2698 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2699 a_n17034_n701# isource_0/VM8D isource_0/VM14D cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X2700 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2701 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2702 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2703 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2704 a_n18150_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2705 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2706 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2707 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2708 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2709 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2710 eigth_mirror_0/I_In eigth_mirror_0/I_In a_n11400_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2711 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2712 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2713 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2714 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2715 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2716 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2717 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2718 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2719 tia_core_0/Out_2 cmirror_channel_0/VN cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2720 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2721 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2722 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2723 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2724 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2725 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2726 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2727 outd_0/InputRef tia_core_0/VM39D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2728 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2729 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2730 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2731 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2732 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2733 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2734 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2735 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2736 cmirror_channel_0/VN cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM6D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2737 cmirror_channel_0/VP outd_0/OutputP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2738 a_n16800_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2739 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2740 a_n22200_n11957# eigth_mirror_0/I_In eigth_mirror_0/I_out_7 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2741 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2742 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2743 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2744 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2745 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2746 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2747 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2748 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2749 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2750 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2751 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2752 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2753 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2754 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2755 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2756 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2757 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2758 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2759 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2760 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2761 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2762 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2763 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2764 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2765 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2766 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2767 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2768 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2769 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2770 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2771 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2772 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X2773 cmirror_channel_0/VP outd_0/OutputN cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2774 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2775 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2776 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2777 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2778 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2779 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2780 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2781 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2782 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2783 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2784 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2785 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2786 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2787 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2788 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2789 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2790 isource_0/VM2D isource_0/VM9D isource_0/VM9D isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2791 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2792 tia_core_0/Input cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM5D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2793 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2794 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2795 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2796 cmirror_channel_0/VN cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM6D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2797 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2798 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2799 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2800 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2801 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2802 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2803 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2804 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2805 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2806 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2807 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2808 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2809 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2810 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2811 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2812 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2813 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2814 outd_0/InputSignal tia_core_0/Input cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2815 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2816 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2817 cmirror_channel_0/VP isource_0/VM8D a_n17034_6079# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2818 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2819 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2820 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2821 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2822 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2823 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2824 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2825 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2826 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2827 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2828 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X2829 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2830 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2831 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2832 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2833 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2834 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2835 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2836 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2837 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2838 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2839 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2840 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2841 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2842 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2843 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2844 cmirror_channel_0/VN a_n15934_n3852# cmirror_channel_0/VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X2845 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2846 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2847 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2848 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2849 a_n12750_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2850 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2851 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2852 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2853 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2854 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2855 cmirror_channel_0/VP a_n5450_n3434# a_n5250_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2856 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2857 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2858 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2859 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2860 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2861 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2862 cmirror_channel_0/VP eigth_mirror_0/I_In a_n19500_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2863 tia_core_0/Out_2 outd_0/InputSignal tia_core_0/Input tia_core_0/Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2864 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2865 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2866 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2867 outd_0/OutputN cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2868 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2869 tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__cap_var_lvt pd=0u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X2870 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2871 outd_0/V_da1_P outd_0/InputSignal outd_0/outd_stage1_0/isource_out outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2872 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2873 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2874 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2875 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2876 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2877 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2878 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2879 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2880 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2881 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2882 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2883 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2884 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2885 cmirror_channel_0/TIA_I_Bias1 a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2886 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2887 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2888 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2889 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2890 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2891 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2892 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2893 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2894 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2895 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2896 isource_0/VM12G a_n22784_2458# cmirror_channel_0/VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X2897 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2898 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2899 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2900 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2901 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2902 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2903 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2904 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2905 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2906 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2907 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2908 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2909 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2910 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2911 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2912 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2913 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2914 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2915 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2916 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2917 tia_core_0/VM36D cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2918 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2919 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2920 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2921 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2922 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2923 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2924 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2925 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2926 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2927 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2928 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2929 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2930 outd_0/InputSignal tia_core_0/Input cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2931 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2932 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2933 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2934 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2935 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2936 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2937 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2938 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2939 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2940 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2941 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2942 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2943 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2944 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2945 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2946 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2947 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2948 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2949 cmirror_channel_0/A_Out_I_Bias a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2950 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2951 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2952 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2953 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2954 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2955 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2956 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2957 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2958 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X2959 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2960 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2961 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2962 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2963 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2964 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2965 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2966 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2967 isource_0/VM2D isource_0/VM2D cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X2968 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2969 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2970 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2971 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2972 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2973 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2974 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2975 cmirror_channel_0/VN tia_core_0/Disable_TIA cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2976 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2977 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2978 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2979 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2980 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2981 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2982 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2983 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2984 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2985 tia_core_0/Out_2 outd_0/InputSignal tia_core_0/Input tia_core_0/Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X2986 outd_0/OutputN cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2987 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2988 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2989 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2990 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2991 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2992 tia_core_0/Input cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM5D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2993 cmirror_channel_0/VP isource_0/VM8D a_n17034_n2971# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2994 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2995 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2996 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2997 outd_0/OutputP cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2998 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2999 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3000 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3001 outd_0/InputRef tia_core_0/VM39D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3002 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3003 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3004 cmirror_channel_0/VN isource_0/VM2D isource_0/VM2D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3005 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3006 tia_core_0/VM5D cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3007 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3008 cmirror_channel_0/VP eigth_mirror_0/I_In a_n22200_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3009 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3010 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3011 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3012 cmirror_channel_0/TIA_I_Bias1 a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3013 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3014 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3015 cmirror_channel_0/VP cmirror_channel_0/VN tia_core_0/Out_2 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3016 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3017 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3018 a_n16800_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3019 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3020 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3021 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3022 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3023 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3024 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3025 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3026 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3027 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3028 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3029 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3030 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3031 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3032 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3033 cmirror_channel_0/VP eigth_mirror_0/I_In a_n20850_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3034 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3035 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3036 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3037 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3038 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3039 cmirror_channel_0/VP isource_0/VM14D isource_0/VM12G isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3040 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3041 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3042 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3043 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3044 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3045 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3046 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3047 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3048 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3049 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3050 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3051 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3052 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3053 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3054 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3055 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3056 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3057 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3058 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3059 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3060 outd_0/outd_stage1_0/isource_out outd_0/InputRef outd_0/V_da1_N outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3061 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3062 a_n4672_n5100# cmirror_channel_0/I_in_channel cmirror_channel_0/TIA_I_Bias2 cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3063 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3064 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3065 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3066 tia_core_0/VM39D outd_0/InputRef tia_core_0/VM31D tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3067 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3068 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3069 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3070 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3071 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3072 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3073 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3074 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3075 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3076 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3077 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3078 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3079 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3080 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3081 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3082 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3083 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3084 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3085 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3086 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3087 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3088 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3089 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3090 isource_0/VM9D isource_0/VM9D isource_0/VM2D isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3091 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3092 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3093 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3094 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3095 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3096 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3097 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3098 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3099 a_n18150_n11957# eigth_mirror_0/I_In eigth_mirror_0/I_out_4 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3100 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3101 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3102 cmirror_channel_0/A_Out_I_Bias a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3103 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3104 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3105 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3106 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3107 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3108 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3109 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3110 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3111 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3112 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3113 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3114 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3115 cmirror_channel_0/VP cmirror_channel_0/VN tia_core_0/Out_2 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3116 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3117 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3118 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3119 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3120 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3121 cmirror_channel_0/VP eigth_mirror_0/I_In a_n11400_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3122 outd_0/OutputP cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3123 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3124 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3125 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3126 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3127 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3128 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3129 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3130 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3131 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3132 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3133 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3134 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3135 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3136 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3137 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3138 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3139 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3140 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3141 a_n19500_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3142 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17268_7820# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3143 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3144 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3145 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3146 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3147 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3148 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3149 isource_0/VM22D a_n35954_n3878# isource_0/VM3D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3150 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3151 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3152 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3153 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3154 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3155 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3156 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3157 isource_0/VM2D isource_0/VM2D cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3158 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3159 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3160 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3161 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3162 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3163 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3164 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3165 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3166 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3167 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3168 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3169 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3170 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3171 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3172 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3173 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3174 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3175 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3176 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3177 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3178 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3179 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3180 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3181 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3182 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3183 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3184 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3185 cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM6D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3186 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3187 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3188 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3189 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3190 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3191 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3192 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3193 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3194 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3195 outd_0/outd_stage1_0/isource_out outd_0/InputSignal outd_0/V_da1_P outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3196 tia_core_0/VM6D cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3197 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3198 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3199 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3200 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3201 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3202 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3203 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3204 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3205 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3206 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3207 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3208 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3209 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3210 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3211 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3212 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3213 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3214 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3215 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3216 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3217 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3218 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3219 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3220 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3221 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3222 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3223 cmirror_channel_0/A_Out_I_Bias a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3224 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3225 isource_0/VM12G isource_0/VM14D cmirror_channel_0/VP isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3226 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3227 a_n18994_26# a_n18464_2458# cmirror_channel_0/VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X3228 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3229 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3230 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3231 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3232 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3233 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3234 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3235 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3236 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3237 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3238 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3239 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3240 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3241 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3242 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3243 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3244 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3245 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3246 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3247 cmirror_channel_0/VN cmirror_channel_0/I_in_channel a_n5512_n5100# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3248 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3249 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3250 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3251 cmirror_channel_0/I_in_channel eigth_mirror_0/I_In a_n12750_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3252 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3253 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3254 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3255 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3256 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3257 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3258 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3259 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3260 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3261 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3262 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3263 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3264 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3265 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3266 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3267 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3268 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3269 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3270 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3271 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3272 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3273 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3274 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3275 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3276 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3277 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3278 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3279 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3280 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3281 a_n17034_n2971# isource_0/VM8D isource_0/VM22D cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X3282 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3283 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3284 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3285 eigth_mirror_0/I_In eigth_mirror_0/I_In a_n11400_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3286 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3287 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3288 cmirror_channel_0/VP isource_0/VM8D sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X3289 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3290 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3291 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3292 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3293 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3294 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3295 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3296 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3297 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3298 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3299 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3300 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3301 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3302 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3303 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3304 tia_core_0/VM36D cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3305 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3306 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3307 a_n11400_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3308 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3309 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3310 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3311 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3312 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3313 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3314 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3315 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3316 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3317 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3318 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3319 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3320 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3321 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3322 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3323 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3324 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3325 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3326 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3327 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3328 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3329 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3330 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3331 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3332 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3333 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3334 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3335 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3336 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3337 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3338 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3339 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3340 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3341 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3342 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3343 outd_0/InputRef tia_core_0/VM39D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3344 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3345 tia_core_0/VM36D cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM39D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3346 a_n12750_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3347 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3348 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3349 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3350 cmirror_channel_0/VP outd_0/OutputN cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3351 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3352 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3353 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3354 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3355 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3356 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3357 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3358 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3359 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3360 isource_0/VM2D isource_0/VM2D cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3361 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3362 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3363 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3364 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3365 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3366 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3367 a_n4672_n5100# cmirror_channel_0/I_in_channel cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3368 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3369 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3370 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3371 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3372 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3373 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3374 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3375 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3376 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3377 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3378 cmirror_channel_0/VP eigth_mirror_0/I_In a_n16800_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3379 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3380 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3381 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3382 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3383 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3384 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3385 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3386 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3387 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3388 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3389 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3390 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3391 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3392 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3393 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3394 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3395 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3396 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3397 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3398 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3399 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3400 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3401 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3402 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3403 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3404 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3405 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3406 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3407 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3408 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3409 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3410 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3411 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3412 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3413 cmirror_channel_0/VN cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM5D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3414 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3415 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3416 eigth_mirror_0/I_In isource_0/VM22D a_n35954_n3878# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3417 cmirror_channel_0/VP eigth_mirror_0/I_In a_n18150_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3418 isource_0/VM2D isource_0/VM9D isource_0/VM9D isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3419 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3420 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3421 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3422 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3423 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3424 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3425 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3426 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3427 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3428 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3429 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3430 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3431 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3432 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3433 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3434 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3435 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3436 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3437 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3438 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3439 outd_0/V_da1_P outd_0/InputSignal outd_0/outd_stage1_0/isource_out outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3440 cmirror_channel_0/VP eigth_mirror_0/I_In a_n14100_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3441 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3442 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3443 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3444 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3445 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3446 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3447 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3448 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3449 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3450 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3451 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3452 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3453 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3454 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3455 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3456 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3457 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3458 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3459 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3460 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3461 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3462 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3463 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3464 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3465 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3466 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3467 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3468 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3469 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3470 isource_0/VM3D a_n35954_n3878# isource_0/VM22D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3471 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3472 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3473 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3474 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3475 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3476 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3477 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3478 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3479 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3480 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3481 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3482 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3483 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3484 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3485 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3486 cmirror_channel_0/VP eigth_mirror_0/I_In a_n20850_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3487 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3488 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3489 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3490 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3491 cmirror_channel_0/VP a_n5450_n3434# a_n5250_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3492 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3493 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3494 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3495 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3496 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3497 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3498 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3499 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3500 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3501 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3502 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3503 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3504 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3505 cmirror_channel_0/TIA_I_Bias1 a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3506 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3507 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3508 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3509 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3510 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3511 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3512 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3513 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3514 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3515 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3516 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3517 isource_0/VM8D isource_0/VM9D isource_0/VM11D isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3518 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3519 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3520 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3521 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3522 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3523 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3524 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3525 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3526 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3527 a_n16800_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3528 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3529 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3530 a_n17034_n701# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3531 a_n17034_n701# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3532 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3533 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3534 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3535 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3536 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3537 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3538 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3539 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3540 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3541 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3542 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3543 isource_0/VM9D isource_0/VM9D isource_0/VM2D isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3544 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3545 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3546 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3547 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3548 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3549 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3550 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3551 outd_0/outd_stage1_0/isource_out outd_0/InputRef outd_0/V_da1_N outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3552 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3553 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3554 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3555 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3556 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3557 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3558 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3559 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3560 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3561 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3562 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3563 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3564 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3565 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3566 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3567 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3568 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3569 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3570 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3571 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3572 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3573 cmirror_channel_0/TIA_I_Bias1 tia_core_0/Disable_TIA cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3574 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3575 a_n21114_26# a_n20584_2458# cmirror_channel_0/VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X3576 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3577 isource_0/VM8D a_n25012_12290# cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X3578 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3579 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3580 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3581 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3582 outd_0/V_da2_N cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3583 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3584 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3585 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3586 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3587 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3588 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3589 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3590 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3591 a_n11400_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3592 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3593 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3594 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3595 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3596 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3597 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3598 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3599 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3600 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3601 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3602 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3603 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3604 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3605 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3606 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3607 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3608 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3609 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3610 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3611 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3612 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3613 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3614 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3615 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3616 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3617 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3618 outd_0/OutputN cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3619 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3620 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3621 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3622 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3623 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3624 outd_0/outd_stage1_0/isource_out outd_0/InputRef outd_0/V_da1_N outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3625 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3626 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3627 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3628 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3629 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3630 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3631 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3632 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3633 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3634 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3635 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3636 cmirror_channel_0/VN cmirror_channel_0/VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3637 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3638 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3639 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3640 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3641 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3642 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3643 a_n17034_n2971# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3644 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3645 tia_core_0/VM5D cmirror_channel_0/TIA_I_Bias1 tia_core_0/Input cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3646 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3647 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3648 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3649 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3650 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3651 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3652 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3653 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3654 a_n19500_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3655 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3656 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3657 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3658 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3659 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3660 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3661 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3662 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3663 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3664 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3665 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3666 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3667 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3668 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3669 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3670 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3671 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3672 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3673 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3674 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3675 a_n12750_n11957# eigth_mirror_0/I_In cmirror_channel_0/I_in_channel cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3676 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3677 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3678 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3679 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3680 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3681 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3682 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3683 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3684 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3685 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3686 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3687 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3688 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3689 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3690 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3691 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3692 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3693 outd_0/OutputP cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3694 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3695 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3696 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3697 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3698 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3699 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3700 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3701 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3702 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3703 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3704 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3705 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3706 a_n17034_n701# isource_0/VM8D isource_0/VM14D cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X3707 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3708 a_n11400_n11957# eigth_mirror_0/I_In eigth_mirror_0/I_In cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3709 cmirror_channel_0/VP eigth_mirror_0/I_In a_n19500_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3710 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3711 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3712 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3713 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3714 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3715 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3716 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3717 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3718 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3719 a_n14100_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3720 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3721 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3722 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3723 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3724 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3725 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3726 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3727 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3728 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3729 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3730 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3731 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3732 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3733 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3734 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3735 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3736 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3737 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3738 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3739 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3740 tia_core_0/VM31D outd_0/InputRef tia_core_0/VM39D tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3741 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3742 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3743 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3744 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3745 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3746 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3747 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3748 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3749 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3750 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3751 a_n17034_6079# isource_0/VM8D isource_0/VM8D cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X3752 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3753 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3754 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3755 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3756 cmirror_channel_0/VP cmirror_channel_0/VN tia_core_0/VM31D cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3757 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3758 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3759 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3760 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3761 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3762 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3763 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3764 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3765 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3766 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3767 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3768 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3769 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3770 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3771 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3772 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3773 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3774 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3775 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3776 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3777 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3778 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3779 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3780 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3781 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3782 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3783 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3784 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3785 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3786 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3787 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3788 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3789 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3790 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3791 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3792 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3793 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3794 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3795 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3796 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3797 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3798 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3799 tia_core_0/Input outd_0/InputSignal tia_core_0/Out_2 tia_core_0/Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3800 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3801 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3802 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3803 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3804 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3805 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3806 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3807 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3808 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3809 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3810 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3811 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3812 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3813 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3814 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3815 a_17268_7820# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3816 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3817 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3818 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3819 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3820 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3821 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3822 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3823 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3824 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3825 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3826 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3827 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3828 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3829 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3830 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3831 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3832 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3833 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3834 cmirror_channel_0/VP eigth_mirror_0/I_In a_n16800_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3835 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3836 a_n19500_n11957# eigth_mirror_0/I_In eigth_mirror_0/I_out_5 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3837 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3838 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3839 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3840 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3841 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3842 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3843 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3844 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3845 cmirror_channel_0/VN isource_0/VM2D isource_0/VM2D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3846 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3847 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3848 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3849 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3850 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3851 a_n20850_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3852 isource_0/VM2D isource_0/VM9D isource_0/VM9D isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3853 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3854 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3855 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3856 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3857 cmirror_channel_0/VP eigth_mirror_0/I_In a_n15450_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3858 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3859 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3860 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3861 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3862 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3863 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3864 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3865 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3866 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3867 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3868 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3869 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3870 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3871 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3872 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3873 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3874 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3875 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3876 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3877 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3878 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3879 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3880 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3881 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3882 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3883 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3884 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3885 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3886 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3887 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3888 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3889 outd_0/V_da1_N outd_0/InputRef outd_0/outd_stage1_0/isource_out outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3890 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3891 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3892 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3893 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3894 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3895 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3896 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3897 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3898 tia_core_0/Input outd_0/InputSignal tia_core_0/Out_2 tia_core_0/Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3899 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3900 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3901 cmirror_channel_0/VP isource_0/VM8D a_n17034_6079# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3902 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3903 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3904 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3905 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3906 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3907 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3908 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3909 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3910 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3911 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3912 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3913 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3914 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3915 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3916 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3917 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3918 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3919 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3920 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3921 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3922 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3923 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3924 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3925 cmirror_channel_0/VP outd_0/V_da2_N cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3926 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3927 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3928 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3929 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3930 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3931 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3932 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3933 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3934 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3935 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3936 outd_0/InputRef tia_core_0/VM39D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3937 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3938 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3939 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3940 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3941 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3942 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3943 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3944 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3945 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3946 cmirror_channel_0/VP eigth_mirror_0/I_In a_n11400_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3947 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3948 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3949 a_n19500_n11957# eigth_mirror_0/I_In eigth_mirror_0/I_out_5 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3950 cmirror_channel_0/VP isource_0/VM8D a_n17034_n2971# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3951 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3952 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3953 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3954 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3955 a_n5450_n3434# a_n5450_n3434# a_n5250_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3956 isource_0/VM8D isource_0/VM9D isource_0/VM11D isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3957 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3958 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3959 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3960 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3961 tia_core_0/VM31D outd_0/InputRef tia_core_0/VM39D tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3962 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3963 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3964 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3965 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3966 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3967 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3968 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3969 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3970 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3971 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3972 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3973 cmirror_channel_0/VP eigth_mirror_0/I_In a_n20850_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3974 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3975 cmirror_channel_0/VP eigth_mirror_0/I_In a_n12750_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3976 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3977 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3978 cmirror_channel_0/VP a_n5450_n3434# a_n5250_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3979 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3980 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3981 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3982 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3983 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3984 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3985 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3986 outd_0/InputSignal tia_core_0/Input cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3987 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3988 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3989 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3990 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3991 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3992 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3993 tia_core_0/VM39D cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM36D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3994 eigth_mirror_0/I_In isource_0/VM22D a_n35954_n3878# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3995 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3996 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3997 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3998 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3999 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4000 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4001 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4002 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4003 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4004 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4005 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4006 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4007 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4008 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4009 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4010 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4011 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4012 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4013 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4014 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4015 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4016 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4017 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4018 cmirror_channel_0/VN isource_0/VM2D isource_0/VM2D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4019 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4020 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4021 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4022 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4023 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4024 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4025 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4026 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4027 tia_core_0/VM39D outd_0/InputRef tia_core_0/VM31D tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4028 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4029 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4030 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4031 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4032 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4033 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4034 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4035 cmirror_channel_0/VN cmirror_channel_0/VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4036 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4037 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4038 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4039 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4040 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4041 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4042 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4043 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4044 a_n35954_n3878# isource_0/VM22D eigth_mirror_0/I_In cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4045 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4046 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4047 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4048 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4049 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4050 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4051 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4052 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4053 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4054 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4055 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4056 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4057 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4058 cmirror_channel_0/VN isource_0/VM2D isource_0/VM2D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4059 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4060 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4061 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4062 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4063 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4064 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4065 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4066 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4067 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4068 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4069 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4070 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4071 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4072 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4073 a_n5450_n3434# a_n5450_n3434# a_n5250_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4074 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4075 a_n11400_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4076 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4077 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4078 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4079 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4080 a_n17034_n701# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4081 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4082 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4083 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4084 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4085 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4086 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4087 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4088 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4089 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4090 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4091 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4092 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4093 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4094 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4095 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4096 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4097 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4098 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4099 outd_0/InputSignal tia_core_0/Input cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4100 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4101 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4102 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4103 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4104 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4105 a_n5512_n5100# cmirror_channel_0/I_in_channel cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4106 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4107 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4108 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4109 tia_core_0/VM39D outd_0/InputRef tia_core_0/VM31D tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4110 outd_0/InputSignal tia_core_0/Input cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4111 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4112 a_n4672_n5100# cmirror_channel_0/I_in_channel cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4113 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4114 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4115 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4116 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4117 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4118 outd_0/OutputP cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4119 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4120 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4121 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4122 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4123 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4124 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4125 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4126 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4127 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4128 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4129 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4130 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4131 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4132 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4133 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4134 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4135 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4136 isource_0/VM9D isource_0/VM9D isource_0/VM2D isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4137 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4138 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4139 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4140 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4141 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4142 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4143 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4144 cmirror_channel_0/VN cmirror_channel_0/I_in_channel sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4145 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4146 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4147 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4148 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4149 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4150 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4151 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4152 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4153 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4154 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4155 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4156 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4157 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4158 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4159 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4160 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4161 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4162 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4163 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4164 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4165 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4166 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4167 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4168 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4169 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4170 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4171 outd_0/OutputN cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4172 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4173 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4174 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4175 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4176 outd_0/InputRef tia_core_0/VM39D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4177 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4178 tia_core_0/VM36D cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM39D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4179 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4180 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4181 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4182 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4183 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4184 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4185 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4186 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4187 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4188 a_n22200_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4189 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4190 isource_0/VM12G isource_0/VM14D cmirror_channel_0/VP isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4191 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4192 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4193 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4194 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4195 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4196 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4197 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4198 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4199 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4200 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4201 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4202 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4203 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4204 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4205 a_n14100_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4206 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4207 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4208 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4209 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4210 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4211 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4212 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4213 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4214 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4215 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4216 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4217 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4218 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4219 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4220 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4221 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4222 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4223 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4224 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4225 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4226 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4227 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4228 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4229 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4230 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4231 outd_0/InputSignal tia_core_0/Input cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4232 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4233 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4234 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4235 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4236 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4237 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4238 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4239 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4240 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4241 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4242 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4243 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4244 cmirror_channel_0/VP eigth_mirror_0/I_In a_n18150_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4245 a_n35954_n3878# isource_0/VM22D eigth_mirror_0/I_In cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4246 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4247 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4248 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4249 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4250 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4251 cmirror_channel_0/VN isource_0/VM2D isource_0/VM2D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4252 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4253 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4254 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4255 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4256 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4257 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4258 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4259 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4260 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4261 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4262 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4263 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4264 outd_0/OutputP cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4265 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4266 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4267 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4268 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4269 cmirror_channel_0/VP eigth_mirror_0/I_In a_n14100_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4270 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4271 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4272 eigth_mirror_0/I_out_6 eigth_mirror_0/I_In a_n20850_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4273 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4274 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4275 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4276 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4277 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4278 tia_core_0/VM6D cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4279 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4280 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4281 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4282 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4283 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4284 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4285 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4286 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4287 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4288 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4289 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4290 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4291 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4292 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4293 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4294 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4295 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4296 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4297 outd_0/OutputP cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4298 cmirror_channel_0/VP eigth_mirror_0/I_In a_n12750_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4299 tia_core_0/VM6D cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4300 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4301 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4302 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4303 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4304 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4305 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4306 tia_core_0/Out_2 outd_0/InputSignal tia_core_0/Input tia_core_0/Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4307 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4308 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4309 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4310 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4311 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4312 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4313 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4314 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4315 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4316 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4317 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4318 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4319 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4320 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4321 cmirror_channel_0/A_Out_I_Bias a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4322 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4323 outd_0/InputRef tia_core_0/VM39D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4324 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4325 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4326 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4327 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4328 cmirror_channel_0/VP eigth_mirror_0/I_In a_n16800_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4329 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4330 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4331 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4332 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4333 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4334 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4335 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4336 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4337 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4338 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4339 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4340 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4341 isource_0/VM8D isource_0/VM9D isource_0/VM11D isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4342 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4343 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4344 tia_core_0/VM39D outd_0/InputRef tia_core_0/VM31D tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4345 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4346 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4347 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4348 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4349 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4350 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4351 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4352 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4353 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4354 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4355 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4356 cmirror_channel_0/VP eigth_mirror_0/I_In a_n15450_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4357 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4358 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4359 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4360 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4361 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4362 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4363 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4364 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4365 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4366 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4367 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4368 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4369 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4370 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4371 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4372 cmirror_channel_0/VP isource_0/VM14D isource_0/VM12G isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4373 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4374 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4375 tia_core_0/VM31D cmirror_channel_0/VN cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4376 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4377 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4378 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4379 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4380 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4381 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4382 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4383 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4384 cmirror_channel_0/VP cmirror_channel_0/VN tia_core_0/VM31D cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4385 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4386 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4387 a_n14100_n11957# eigth_mirror_0/I_In eigth_mirror_0/I_out_1 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4388 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4389 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4390 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4391 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4392 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4393 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4394 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4395 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4396 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4397 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4398 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4399 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4400 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4401 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4402 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4403 cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4404 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4405 cmirror_channel_0/VP outd_0/V_da2_N cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4406 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4407 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4408 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4409 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4410 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4411 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4412 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4413 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4414 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4415 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4416 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4417 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4418 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4419 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4420 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4421 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4422 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4423 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4424 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4425 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4426 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4427 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4428 outd_0/V_da1_N outd_0/InputRef outd_0/outd_stage1_0/isource_out outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4429 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4430 cmirror_channel_0/VN cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM6D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4431 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4432 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4433 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4434 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4435 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4436 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4437 a_n17034_8339# isource_0/VM8D isource_0/VM9D cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X4438 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4439 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4440 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4441 isource_0/VM2D isource_0/VM9D isource_0/VM9D isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4442 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4443 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4444 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4445 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4446 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4447 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4448 cmirror_channel_0/VP isource_0/VM8D a_n17034_6079# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4449 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4450 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4451 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4452 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4453 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4454 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4455 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4456 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4457 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4458 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4459 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4460 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4461 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4462 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4463 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4464 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4465 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4466 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4467 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4468 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4469 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4470 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4471 cmirror_channel_0/A_Out_I_Bias a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4472 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4473 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4474 cmirror_channel_0/VN cmirror_channel_0/VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4475 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4476 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4477 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4478 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4479 cmirror_channel_0/TIA_I_Bias1 a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4480 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4481 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4482 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4483 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4484 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4485 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4486 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4487 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4488 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4489 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4490 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4491 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4492 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4493 a_n17034_n701# isource_0/VM8D isource_0/VM14D cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X4494 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4495 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4496 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4497 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4498 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4499 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4500 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4501 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4502 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4503 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4504 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4505 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4506 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4507 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4508 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4509 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4510 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4511 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4512 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4513 isource_0/VM3D a_n35954_n3878# isource_0/VM22D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4514 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4515 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4516 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4517 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4518 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4519 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4520 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4521 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4522 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4523 a_n5512_n5100# cmirror_channel_0/I_in_channel a_n5450_n3434# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4524 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4525 isource_0/VM2D isource_0/VM9D isource_0/VM9D isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4526 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4527 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4528 outd_0/V_da1_P cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
X4529 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4530 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4531 a_n18150_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4532 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4533 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4534 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4535 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4536 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4537 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4538 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4539 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4540 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4541 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4542 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4543 tia_core_0/Input outd_0/InputSignal tia_core_0/Out_2 tia_core_0/Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4544 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4545 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4546 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4547 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4548 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4549 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4550 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4551 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4552 outd_0/V_da1_N cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
X4553 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4554 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4555 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4556 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4557 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4558 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4559 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4560 outd_0/V_da1_P cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
X4561 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4562 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4563 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4564 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4565 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4566 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4567 cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/A_Out_I_Bias a_17268_7820# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4568 isource_0/VM3D isource_0/VM3G cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4569 a_n25012_12290# isource_0/VM11D cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X4570 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4571 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4572 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4573 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4574 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4575 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4576 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4577 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4578 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4579 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4580 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4581 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4582 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4583 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4584 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4585 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4586 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4587 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4588 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4589 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4590 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4591 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4592 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4593 cmirror_channel_0/A_Out_I_Bias a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4594 a_n17034_n701# isource_0/VM8D isource_0/VM14D cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X4595 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4596 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4597 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4598 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4599 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4600 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4601 outd_0/OutputN cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4602 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4603 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4604 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4605 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4606 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4607 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4608 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4609 cmirror_channel_0/TIA_I_Bias1 a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4610 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4611 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4612 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4613 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4614 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4615 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4616 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4617 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4618 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4619 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4620 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4621 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4622 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4623 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4624 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4625 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4626 cmirror_channel_0/VP isource_0/VM8D a_n17034_8339# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4627 a_n17034_6079# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4628 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4629 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4630 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4631 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4632 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4633 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4634 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4635 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4636 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4637 a_n17034_n701# isource_0/VM8D isource_0/VM14D cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X4638 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4639 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4640 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4641 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4642 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4643 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4644 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4645 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4646 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4647 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4648 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4649 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4650 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4651 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4652 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4653 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4654 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4655 eigth_mirror_0/I_out_2 eigth_mirror_0/I_In a_n15450_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4656 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4657 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4658 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4659 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4660 cmirror_channel_0/VP a_n5450_n3434# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4661 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4662 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4663 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4664 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4665 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4666 isource_0/VM2D isource_0/VM2D cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4667 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4668 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4669 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4670 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4671 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4672 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4673 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4674 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4675 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4676 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4677 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4678 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4679 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4680 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4681 a_n17034_n701# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4682 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4683 cmirror_channel_0/VN cmirror_channel_0/I_in_channel a_n4672_n5100# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4684 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4685 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4686 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4687 cmirror_channel_0/VP eigth_mirror_0/I_In a_n15450_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4688 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4689 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4690 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4691 a_n5250_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4692 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4693 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4694 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4695 eigth_mirror_0/I_In isource_0/VM22D a_n35954_n3878# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4696 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4697 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4698 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4699 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4700 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4701 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4702 a_n25012_12290# isource_0/VM11D cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X4703 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4704 outd_0/V_da2_P cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4705 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4706 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4707 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4708 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4709 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4710 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4711 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4712 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4713 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4714 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4715 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4716 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4717 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4718 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4719 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4720 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4721 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4722 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4723 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4724 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4725 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4726 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4727 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4728 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4729 tia_core_0/Input outd_0/InputSignal tia_core_0/Out_2 tia_core_0/Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4730 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4731 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4732 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4733 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4734 isource_0/VM11D isource_0/VM9D isource_0/VM8D isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4735 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4736 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4737 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4738 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4739 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4740 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4741 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4742 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4743 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4744 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4745 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4746 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4747 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4748 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4749 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4750 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4751 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4752 outd_0/OutputN cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4753 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4754 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4755 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4756 cmirror_channel_0/A_Out_I_Bias a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4757 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4758 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4759 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4760 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4761 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4762 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4763 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4764 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4765 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4766 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4767 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4768 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4769 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4770 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4771 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4772 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4773 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4774 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4775 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4776 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4777 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4778 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4779 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4780 cmirror_channel_0/VN isource_0/VM12G isource_0/VM14D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4781 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4782 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4783 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4784 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4785 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4786 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4787 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4788 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4789 outd_0/V_da1_N cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
X4790 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4791 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4792 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4793 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4794 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4795 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4796 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4797 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4798 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4799 outd_0/InputRef tia_core_0/VM39D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4800 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4801 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4802 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4803 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4804 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4805 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4806 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4807 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4808 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4809 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4810 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4811 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4812 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4813 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4814 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4815 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4816 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4817 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4818 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4819 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4820 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4821 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4822 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4823 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4824 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4825 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4826 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4827 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4828 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4829 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4830 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4831 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4832 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4833 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4834 a_n35954_n3878# isource_0/VM22D eigth_mirror_0/I_In cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4835 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4836 cmirror_channel_0/VP a_n5450_n3434# a_n5250_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4837 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4838 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4839 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4840 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4841 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4842 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4843 outd_0/V_da2_P cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4844 eigth_mirror_0/I_out_6 eigth_mirror_0/I_In a_n20850_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4845 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4846 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4847 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4848 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4849 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4850 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4851 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4852 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4853 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4854 isource_0/VM22D a_n35954_n3878# isource_0/VM3D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4855 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4856 a_n5512_n5100# cmirror_channel_0/I_in_channel cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4857 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4858 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4859 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4860 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4861 a_n20850_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4862 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4863 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4864 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4865 outd_0/OutputP cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4866 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4867 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4868 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4869 cmirror_channel_0/A_Out_I_Bias a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4870 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4871 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4872 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4873 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4874 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4875 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4876 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4877 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4878 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4879 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4880 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4881 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4882 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4883 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4884 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4885 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4886 eigth_mirror_0/I_In isource_0/VM22D a_n35954_n3878# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4887 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4888 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4889 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4890 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4891 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4892 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4893 cmirror_channel_0/VP outd_0/OutputN cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4894 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4895 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4896 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4897 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4898 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4899 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4900 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4901 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4902 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4903 isource_0/VM2D isource_0/VM9D isource_0/VM9D isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4904 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4905 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4906 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4907 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4908 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4909 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4910 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4911 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4912 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4913 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4914 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4915 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4916 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4917 isource_0/VM2D isource_0/VM2D cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4918 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4919 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4920 cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM6D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4921 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4922 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4923 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4924 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4925 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4926 outd_0/InputRef tia_core_0/VM39D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4927 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4928 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4929 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4930 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4931 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4932 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4933 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4934 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4935 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4936 cmirror_channel_0/TIA_I_Bias1 a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4937 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4938 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4939 tia_core_0/VM36D cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM39D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4940 a_n12750_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4941 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4942 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4943 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4944 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4945 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4946 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4947 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4948 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4949 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4950 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4951 cmirror_channel_0/VP isource_0/VM14D isource_0/VM12G isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4952 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4953 outd_0/outd_stage1_0/isource_out outd_0/InputRef outd_0/V_da1_N outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4954 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4955 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4956 outd_0/InputSignal tia_core_0/Input cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4957 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4958 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4959 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4960 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4961 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4962 isource_0/VM3G a_n22784_2458# cmirror_channel_0/VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X4963 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4964 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4965 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4966 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4967 a_n17034_n701# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4968 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4969 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4970 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4971 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4972 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4973 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4974 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4975 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4976 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4977 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4978 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4979 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4980 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4981 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4982 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4983 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4984 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4985 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4986 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4987 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4988 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4989 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4990 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4991 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4992 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4993 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4994 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4995 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4996 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4997 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4998 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4999 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5000 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5001 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5002 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5003 cmirror_channel_0/VP eigth_mirror_0/I_In a_n22200_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5004 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5005 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5006 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5007 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5008 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5009 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5010 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5011 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5012 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5013 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5014 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5015 a_n35954_n3878# isource_0/VM22D eigth_mirror_0/I_In cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5016 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5017 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5018 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5019 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5020 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5021 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5022 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5023 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5024 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5025 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5026 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5027 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5028 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5029 cmirror_channel_0/TIA_I_Bias1 a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5030 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5031 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5032 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5033 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5034 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5035 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5036 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5037 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5038 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5039 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5040 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5041 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5042 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5043 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5044 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5045 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5046 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5047 outd_0/InputSignal tia_core_0/Input cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5048 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5049 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5050 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5051 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5052 tia_core_0/Out_2 outd_0/InputSignal tia_core_0/Input tia_core_0/Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5053 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5054 eigth_mirror_0/I_In isource_0/VM22D a_n35954_n3878# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5055 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5056 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5057 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5058 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5059 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5060 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5061 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5062 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5063 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5064 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5065 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5066 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5067 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5068 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5069 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5070 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5071 a_n16800_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5072 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5073 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5074 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5075 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5076 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5077 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5078 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5079 a_n17034_8339# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5080 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5081 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5082 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5083 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5084 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5085 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5086 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5087 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5088 a_n12750_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5089 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5090 cmirror_channel_0/VN cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM36D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5091 isource_0/VM11D isource_0/VM9D isource_0/VM8D isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5092 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5093 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5094 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5095 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5096 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5097 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5098 cmirror_channel_0/A_Out_I_Bias a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5099 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5100 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5101 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5102 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5103 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5104 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5105 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5106 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5107 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5108 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5109 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5110 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5111 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5112 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5113 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5114 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5115 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5116 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5117 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5118 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5119 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5120 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5121 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5122 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5123 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5124 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5125 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5126 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5127 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5128 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5129 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5130 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5131 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5132 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5133 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5134 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5135 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5136 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5137 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5138 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5139 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5140 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5141 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5142 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5143 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5144 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5145 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5146 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5147 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5148 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5149 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5150 tia_core_0/VM31D outd_0/InputRef tia_core_0/VM39D tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5151 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5152 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5153 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5154 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5155 outd_0/OutputN cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5156 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5157 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5158 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5159 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5160 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5161 a_n17034_n701# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5162 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5163 cmirror_channel_0/VP eigth_mirror_0/I_In a_n15450_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5164 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5165 outd_0/V_da1_N outd_0/InputRef outd_0/outd_stage1_0/isource_out outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5166 a_n5250_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5167 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5168 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5169 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5170 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5171 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5172 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5173 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5174 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5175 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5176 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5177 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5178 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5179 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5180 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5181 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5182 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5183 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5184 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5185 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5186 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5187 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5188 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5189 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5190 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5191 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5192 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5193 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5194 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5195 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5196 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5197 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5198 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5199 eigth_mirror_0/I_out_2 eigth_mirror_0/I_In a_n15450_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5200 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5201 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5202 a_n19500_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5203 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5204 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5205 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5206 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5207 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5208 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5209 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5210 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5211 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5212 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5213 cmirror_channel_0/A_Out_I_Bias a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5214 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5215 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5216 a_n15450_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5217 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5218 a_n20850_n11957# eigth_mirror_0/I_In eigth_mirror_0/I_out_6 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5219 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5220 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5221 a_n17034_n701# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5222 a_n17034_n701# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5223 a_n5250_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5224 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5225 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5226 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5227 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5228 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5229 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5230 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5231 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5232 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5233 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5234 cmirror_channel_0/VN isource_0/VM3G isource_0/VM3D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X5235 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5236 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5237 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5238 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5239 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5240 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5241 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5242 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5243 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5244 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5245 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5246 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5247 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5248 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5249 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5250 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5251 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5252 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5253 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5254 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5255 a_n17034_n701# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5256 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5257 cmirror_channel_0/TIA_I_Bias1 a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5258 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5259 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5260 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5261 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5262 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5263 a_n22200_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5264 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5265 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5266 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5267 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5268 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5269 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5270 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5271 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5272 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5273 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5274 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5275 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5276 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5277 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5278 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5279 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5280 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5281 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5282 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5283 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5284 outd_0/OutputN cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5285 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5286 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5287 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5288 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5289 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5290 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5291 outd_0/OutputP cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5292 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5293 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5294 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5295 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5296 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5297 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5298 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5299 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5300 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5301 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5302 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5303 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5304 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5305 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5306 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5307 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5308 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5309 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5310 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5311 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5312 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5313 cmirror_channel_0/VP isource_0/VM8D a_n17034_8339# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5314 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5315 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5316 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5317 cmirror_channel_0/A_Out_I_Bias a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5318 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5319 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5320 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5321 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5322 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5323 cmirror_channel_0/VN tia_core_0/Disable_TIA cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5324 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5325 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5326 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5327 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5328 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5329 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5330 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5331 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5332 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5333 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5334 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5335 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5336 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5337 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5338 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5339 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5340 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5341 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5342 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5343 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5344 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5345 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5346 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5347 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5348 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5349 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5350 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5351 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5352 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5353 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5354 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5355 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5356 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5357 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5358 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5359 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5360 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5361 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5362 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5363 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5364 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5365 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5366 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5367 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5368 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5369 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5370 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5371 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5372 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5373 outd_0/InputRef tia_core_0/VM39D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5374 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5375 cmirror_channel_0/TIA_I_Bias1 a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5376 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5377 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5378 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5379 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5380 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5381 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5382 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5383 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5384 cmirror_channel_0/VP isource_0/VM14D isource_0/VM12G isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5385 a_n19500_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5386 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5387 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5388 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5389 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5390 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5391 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5392 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5393 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5394 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5395 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5396 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5397 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5398 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5399 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5400 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5401 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5402 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5403 cmirror_channel_0/VN cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM5D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5404 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5405 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5406 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5407 outd_0/InputSignal tia_core_0/Input cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5408 outd_0/OutputP cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5409 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5410 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5411 outd_0/V_da1_P outd_0/InputSignal outd_0/outd_stage1_0/isource_out outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5412 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5413 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5414 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5415 outd_0/InputSignal tia_core_0/Input cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5416 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5417 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5418 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5419 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5420 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5421 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5422 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5423 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5424 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5425 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5426 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5427 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5428 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5429 cmirror_channel_0/A_Out_I_Bias a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5430 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5431 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5432 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5433 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5434 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5435 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5436 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5437 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5438 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5439 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5440 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5441 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5442 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5443 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5444 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5445 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5446 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5447 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5448 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5449 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5450 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5451 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5452 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5453 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5454 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5455 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5456 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5457 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5458 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5459 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5460 a_n17524_n6284# a_n16994_n3852# cmirror_channel_0/VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X5461 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5462 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5463 cmirror_channel_0/VN isource_0/VM12G isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X5464 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5465 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5466 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5467 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5468 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5469 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5470 tia_core_0/VM39D outd_0/InputRef tia_core_0/VM31D tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5471 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5472 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5473 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5474 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5475 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5476 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5477 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5478 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5479 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5480 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5481 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5482 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5483 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5484 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5485 eigth_mirror_0/I_out_3 eigth_mirror_0/I_In a_n16800_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5486 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5487 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5488 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5489 a_n15450_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5490 tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__cap_var_lvt pd=0u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X5491 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5492 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5493 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5494 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5495 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5496 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5497 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5498 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5499 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5500 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5501 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5502 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5503 a_n35954_n3878# isource_0/VM22D eigth_mirror_0/I_In cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5504 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5505 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5506 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5507 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5508 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5509 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5510 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5511 outd_0/InputRef tia_core_0/VM39D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5512 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5513 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5514 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5515 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5516 a_n14100_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5517 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5518 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5519 outd_0/InputSignal tia_core_0/Input cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5520 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5521 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5522 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5523 outd_0/InputSignal tia_core_0/Input cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5524 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5525 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5526 tia_core_0/VM6D cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5527 cmirror_channel_0/VP isource_0/VM8D a_n17034_6079# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5528 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5529 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5530 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5531 cmirror_channel_0/VP eigth_mirror_0/I_In a_n20850_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5532 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5533 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5534 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5535 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5536 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5537 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5538 tia_core_0/VM39D outd_0/InputRef tia_core_0/VM31D tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5539 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5540 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5541 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5542 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5543 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5544 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5545 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5546 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5547 isource_0/VM2D isource_0/VM2D cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X5548 tia_core_0/VM39D cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM36D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5549 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5550 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5551 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5552 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5553 a_n6352_n5100# cmirror_channel_0/I_in_channel cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5554 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5555 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5556 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5557 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5558 isource_0/VM2D isource_0/VM9D isource_0/VM9D isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5559 a_n5512_n5100# cmirror_channel_0/I_in_channel cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5560 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5561 isource_0/VM12G isource_0/VM14D cmirror_channel_0/VP isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5562 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5563 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5564 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5565 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5566 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5567 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5568 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5569 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5570 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5571 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5572 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5573 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5574 cmirror_channel_0/VN isource_0/VM2D isource_0/VM2D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X5575 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5576 cmirror_channel_0/A_Out_I_Bias a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5577 cmirror_channel_0/VN tia_core_0/Disable_TIA tia_core_0/Disable_TIA_B cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=1e+06u
X5578 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5579 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5580 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5581 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5582 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5583 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5584 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5585 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5586 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5587 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5588 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5589 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5590 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5591 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5592 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5593 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5594 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5595 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5596 a_n20054_26# a_n20584_2458# cmirror_channel_0/VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X5597 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5598 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5599 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5600 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5601 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5602 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5603 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5604 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5605 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5606 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5607 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5608 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5609 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5610 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5611 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5612 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5613 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5614 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5615 a_n18150_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5616 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5617 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5618 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5619 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5620 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5621 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5622 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5623 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5624 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5625 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5626 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5627 a_n11400_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5628 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5629 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5630 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5631 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5632 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5633 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5634 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5635 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5636 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5637 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5638 outd_0/InputSignal tia_core_0/Input cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5639 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5640 cmirror_channel_0/VP outd_0/OutputN cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5641 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5642 a_n16800_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5643 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5644 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5645 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5646 outd_0/outd_stage1_0/isource_out outd_0/InputSignal outd_0/V_da1_P outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5647 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5648 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5649 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5650 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5651 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5652 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5653 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5654 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5655 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X5656 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5657 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5658 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5659 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5660 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5661 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5662 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5663 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5664 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5665 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5666 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5667 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5668 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5669 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5670 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5671 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5672 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5673 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5674 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5675 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5676 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5677 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5678 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5679 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5680 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5681 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5682 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5683 a_n17034_6079# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5684 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5685 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5686 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5687 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5688 cmirror_channel_0/A_Out_I_Bias a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5689 cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5690 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5691 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5692 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5693 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5694 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5695 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5696 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5697 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5698 cmirror_channel_0/VP isource_0/VM8D a_n17034_n2971# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5699 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5700 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5701 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5702 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5703 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5704 tia_core_0/VM5D cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5705 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5706 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5707 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5708 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5709 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5710 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5711 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5712 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5713 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5714 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5715 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5716 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5717 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5718 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5719 isource_0/VM2D isource_0/VM2D cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X5720 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5721 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5722 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5723 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5724 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5725 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5726 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5727 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5728 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5729 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5730 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5731 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5732 outd_0/InputRef tia_core_0/VM39D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5733 isource_0/VM12G isource_0/VM14D cmirror_channel_0/VP isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5734 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5735 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5736 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5737 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5738 outd_0/V_da1_N outd_0/InputRef outd_0/outd_stage1_0/isource_out outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5739 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5740 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5741 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5742 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5743 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5744 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5745 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5746 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5747 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5748 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5749 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5750 a_n22200_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5751 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5752 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5753 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5754 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5755 a_n14100_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5756 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5757 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5758 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5759 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5760 cmirror_channel_0/VP eigth_mirror_0/I_In a_n19500_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5761 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5762 tia_core_0/VM5D cmirror_channel_0/TIA_I_Bias1 tia_core_0/Input cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5763 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5764 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5765 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5766 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5767 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5768 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5769 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5770 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5771 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5772 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5773 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5774 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5775 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5776 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5777 cmirror_channel_0/VP tia_core_0/VM40D sky130_fd_pr__cap_mim_m3_2 l=1.8e+07u w=2.5e+07u
X5778 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5779 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5780 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5781 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5782 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5783 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5784 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5785 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5786 a_n17524_n6284# a_n35954_n3878# cmirror_channel_0/VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X5787 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5788 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5789 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5790 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5791 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5792 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5793 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5794 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5795 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5796 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5797 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5798 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5799 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5800 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5801 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5802 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5803 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5804 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5805 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5806 tia_core_0/VM39D outd_0/InputRef tia_core_0/VM31D tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5807 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5808 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5809 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5810 cmirror_channel_0/VP eigth_mirror_0/I_In a_n22200_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5811 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5812 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5813 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5814 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5815 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5816 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5817 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5818 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5819 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5820 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5821 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5822 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5823 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5824 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5825 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5826 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5827 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5828 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5829 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5830 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5831 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5832 cmirror_channel_0/VN cmirror_channel_0/VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5833 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5834 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5835 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5836 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5837 outd_0/OutputP cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5838 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5839 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5840 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5841 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5842 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5843 cmirror_channel_0/VP eigth_mirror_0/I_In a_n20850_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5844 isource_0/VM14D isource_0/VM12G cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X5845 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5846 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5847 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5848 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5849 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5850 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5851 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5852 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5853 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5854 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5855 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5856 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5857 outd_0/V_da2_N cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5858 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5859 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5860 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5861 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5862 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5863 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5864 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5865 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5866 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5867 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5868 cmirror_channel_0/VP outd_0/OutputN cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5869 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5870 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5871 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5872 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5873 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5874 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5875 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5876 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5877 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5878 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5879 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5880 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5881 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5882 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5883 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5884 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5885 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5886 cmirror_channel_0/VN cmirror_channel_0/I_in_channel a_n6352_n5100# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5887 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5888 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5889 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5890 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5891 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5892 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5893 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5894 cmirror_channel_0/VP eigth_mirror_0/I_In a_n16800_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5895 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5896 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5897 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5898 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5899 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5900 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5901 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5902 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5903 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5904 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5905 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5906 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5907 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5908 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5909 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5910 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5911 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5912 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5913 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5914 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5915 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5916 cmirror_channel_0/VP eigth_mirror_0/I_In a_n15450_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5917 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5918 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5919 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5920 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5921 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5922 isource_0/VM2D isource_0/VM9D isource_0/VM9D isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5923 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5924 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5925 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5926 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5927 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5928 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5929 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5930 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5931 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5932 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5933 cmirror_channel_0/VP a_n5450_n3434# a_n5250_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5934 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5935 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5936 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5937 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5938 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5939 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5940 cmirror_channel_0/VP eigth_mirror_0/I_In a_n11400_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5941 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5942 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5943 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5944 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5945 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5946 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5947 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5948 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5949 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5950 cmirror_channel_0/VP isource_0/VM8D a_n17034_n2971# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5951 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5952 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5953 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5954 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5955 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5956 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5957 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5958 isource_0/VM2D isource_0/VM2D cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X5959 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5960 a_n22200_n11957# eigth_mirror_0/I_In eigth_mirror_0/I_out_7 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5961 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5962 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5963 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5964 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5965 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5966 cmirror_channel_0/VP outd_0/V_da2_P cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5967 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5968 cmirror_channel_0/VP outd_0/OutputN cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5969 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5970 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5971 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5972 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5973 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5974 outd_0/V_da1_P outd_0/InputSignal outd_0/outd_stage1_0/isource_out outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5975 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5976 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5977 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5978 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5979 tia_core_0/Input outd_0/InputSignal tia_core_0/Out_2 tia_core_0/Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5980 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5981 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5982 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5983 isource_0/VM22D a_n35954_n3878# isource_0/VM3D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X5984 outd_0/OutputP cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5985 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5986 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5987 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5988 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5989 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5990 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5991 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5992 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5993 a_n6352_n5100# cmirror_channel_0/I_in_channel cmirror_channel_0/I_in_channel cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5994 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5995 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5996 a_n15450_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5997 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5998 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5999 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6000 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6001 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6002 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6003 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6004 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6005 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6006 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6007 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6008 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6009 cmirror_channel_0/VP outd_0/OutputP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X6010 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6011 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6012 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6013 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6014 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6015 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6016 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6017 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6018 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6019 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6020 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6021 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6022 a_n14100_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6023 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6024 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6025 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6026 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6027 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6028 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6029 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6030 tia_core_0/Out_2 cmirror_channel_0/VN cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6031 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6032 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6033 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6034 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6035 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6036 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6037 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6038 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6039 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6040 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6041 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6042 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6043 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6044 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6045 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6046 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6047 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6048 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6049 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6050 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6051 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6052 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6053 eigth_mirror_0/I_out_3 eigth_mirror_0/I_In a_n16800_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6054 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6055 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6056 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6057 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6058 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6059 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6060 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6061 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6062 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6063 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6064 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6065 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6066 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6067 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6068 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6069 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6070 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6071 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6072 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6073 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6074 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6075 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6076 tia_core_0/Input outd_0/InputSignal tia_core_0/Out_2 tia_core_0/Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6077 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6078 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6079 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6080 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6081 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6082 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6083 cmirror_channel_0/VP outd_0/V_da2_P cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X6084 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6085 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6086 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6087 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6088 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6089 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6090 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6091 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6092 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6093 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6094 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6095 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6096 outd_0/InputRef tia_core_0/VM39D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6097 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6098 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6099 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6100 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6101 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6102 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6103 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6104 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6105 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6106 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6107 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6108 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6109 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6110 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6111 cmirror_channel_0/VP outd_0/OutputP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X6112 tia_core_0/VM31D cmirror_channel_0/VN cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6113 a_n18150_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6114 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6115 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6116 tia_core_0/VM31D outd_0/InputRef tia_core_0/VM39D tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6117 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6118 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6119 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6120 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6121 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6122 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6123 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6124 cmirror_channel_0/VN cmirror_channel_0/I_in_channel a_n5512_n5100# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6125 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6126 tia_core_0/Out_2 cmirror_channel_0/VN cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6127 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6128 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6129 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6130 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6131 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6132 a_n16800_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6133 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6134 outd_0/V_da1_P outd_0/InputSignal outd_0/outd_stage1_0/isource_out outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6135 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6136 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6137 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6138 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6139 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6140 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6141 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6142 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6143 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6144 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6145 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6146 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6147 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6148 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6149 outd_0/InputSignal tia_core_0/Input cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6150 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6151 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6152 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6153 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6154 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6155 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6156 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6157 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6158 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6159 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6160 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6161 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6162 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6163 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6164 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6165 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6166 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6167 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6168 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6169 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6170 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6171 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6172 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6173 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6174 cmirror_channel_0/VP eigth_mirror_0/I_In a_n16800_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6175 tia_core_0/VM31D outd_0/InputRef tia_core_0/VM39D tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6176 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6177 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6178 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6179 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6180 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6181 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6182 outd_0/outd_stage1_0/isource_out outd_0/InputSignal outd_0/V_da1_P outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6183 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6184 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6185 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6186 a_n11400_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6187 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6188 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6189 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6190 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6191 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6192 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6193 cmirror_channel_0/VN isource_0/VM11D a_n25012_12290# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X6194 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6195 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6196 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6197 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6198 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6199 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6200 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6201 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6202 cmirror_channel_0/VP eigth_mirror_0/I_In a_n18150_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6203 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6204 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6205 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6206 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6207 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6208 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6209 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6210 a_n17034_n2971# isource_0/VM8D isource_0/VM22D cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X6211 outd_0/outd_stage1_0/isource_out outd_0/InputSignal outd_0/V_da1_P outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6212 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6213 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6214 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6215 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6216 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6217 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6218 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6219 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6220 cmirror_channel_0/VP outd_0/OutputP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X6221 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6222 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6223 cmirror_channel_0/VP isource_0/VM8D a_n17034_8339# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6224 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6225 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6226 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6227 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6228 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6229 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6230 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6231 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6232 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6233 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6234 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6235 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6236 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6237 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6238 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6239 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6240 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6241 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6242 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6243 cmirror_channel_0/VP eigth_mirror_0/I_In a_n19500_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6244 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6245 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6246 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6247 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6248 isource_0/VM8D isource_0/VM9D isource_0/VM11D isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6249 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6250 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6251 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6252 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6253 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6254 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6255 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6256 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6257 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6258 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6259 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6260 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6261 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6262 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6263 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6264 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6265 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6266 isource_0/VM3D a_n35954_n3878# isource_0/VM22D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6267 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6268 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6269 a_n6352_n5100# cmirror_channel_0/I_in_channel cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6270 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6271 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6272 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6273 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6274 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6275 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6276 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6277 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6278 a_n18150_n11957# eigth_mirror_0/I_In eigth_mirror_0/I_out_4 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6279 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6280 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6281 outd_0/V_da1_N outd_0/InputRef outd_0/outd_stage1_0/isource_out outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6282 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6283 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6284 tia_core_0/Out_2 outd_0/InputSignal tia_core_0/Input tia_core_0/Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6285 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6286 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6287 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6288 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6289 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6290 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6291 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6292 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6293 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6294 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6295 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6296 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6297 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6298 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6299 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6300 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6301 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6302 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6303 outd_0/OutputN cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X6304 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6305 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6306 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6307 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6308 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6309 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6310 cmirror_channel_0/VP eigth_mirror_0/I_In a_n14100_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6311 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6312 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6313 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6314 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6315 outd_0/InputRef tia_core_0/VM39D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6316 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6317 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6318 cmirror_channel_0/VN isource_0/VM11D a_n25012_12290# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X6319 outd_0/InputRef tia_core_0/VM39D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6320 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6321 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6322 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6323 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6324 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6325 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6326 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6327 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6328 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6329 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6330 tia_core_0/VM5D cmirror_channel_0/TIA_I_Bias1 tia_core_0/Input cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6331 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6332 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6333 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6334 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6335 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6336 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6337 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6338 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6339 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6340 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6341 tia_core_0/Out_2 outd_0/InputSignal tia_core_0/Input tia_core_0/Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6342 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6343 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6344 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6345 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6346 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6347 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6348 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6349 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6350 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6351 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6352 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6353 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6354 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6355 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6356 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6357 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6358 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6359 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6360 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X6361 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6362 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6363 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6364 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6365 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6366 a_n17034_n701# isource_0/VM8D isource_0/VM14D cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X6367 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6368 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6369 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6370 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6371 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6372 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6373 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6374 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6375 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6376 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6377 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6378 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6379 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6380 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6381 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6382 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6383 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6384 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6385 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6386 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6387 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6388 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6389 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6390 tia_core_0/Input cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM5D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6391 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6392 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6393 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6394 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6395 outd_0/OutputP cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X6396 a_n17034_8339# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6397 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6398 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6399 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6400 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6401 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6402 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6403 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6404 cmirror_channel_0/VP cmirror_channel_0/VN tia_core_0/Out_2 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6405 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6406 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6407 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6408 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6409 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6410 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6411 cmirror_channel_0/VN isource_0/VM2D isource_0/VM2D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6412 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6413 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6414 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6415 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6416 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6417 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6418 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6419 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6420 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6421 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6422 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6423 tia_core_0/Out_2 outd_0/InputSignal tia_core_0/Input tia_core_0/Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6424 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6425 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6426 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6427 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6428 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6429 tia_core_0/VM31D outd_0/InputRef tia_core_0/VM39D tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6430 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6431 isource_0/VM11D isource_0/VM9D isource_0/VM8D isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6432 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6433 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6434 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6435 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6436 cmirror_channel_0/VP outd_0/OutputN cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X6437 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6438 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6439 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6440 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6441 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6442 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6443 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6444 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6445 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6446 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6447 cmirror_channel_0/VN isource_0/VM11D a_n25012_12290# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X6448 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6449 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6450 a_n16800_n11957# eigth_mirror_0/I_In eigth_mirror_0/I_out_3 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6451 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6452 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6453 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6454 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6455 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6456 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6457 a_n17034_n701# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6458 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6459 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6460 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6461 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6462 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6463 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6464 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6465 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6466 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6467 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6468 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6469 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6470 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6471 outd_0/V_da1_P outd_0/InputSignal outd_0/outd_stage1_0/isource_out outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6472 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6473 tia_core_0/Out_2 outd_0/InputSignal tia_core_0/Input tia_core_0/Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6474 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6475 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6476 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6477 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6478 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6479 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6480 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6481 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6482 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6483 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6484 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6485 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6486 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6487 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6488 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6489 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6490 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6491 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6492 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6493 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6494 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6495 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6496 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6497 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6498 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6499 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6500 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6501 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6502 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6503 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6504 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6505 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6506 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6507 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6508 tia_core_0/VM39D outd_0/InputRef tia_core_0/VM31D tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6509 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6510 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6511 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6512 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6513 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6514 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6515 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6516 isource_0/VM8D isource_0/VM9D isource_0/VM11D isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6517 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6518 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6519 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6520 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6521 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6522 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6523 cmirror_channel_0/VN cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM5D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6524 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6525 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6526 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6527 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6528 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6529 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6530 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6531 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6532 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6533 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6534 isource_0/VM12G isource_0/VM14D cmirror_channel_0/VP isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6535 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6536 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6537 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6538 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6539 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6540 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6541 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6542 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6543 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6544 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6545 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6546 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6547 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6548 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6549 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6550 isource_0/VM12D isource_0/VM12G cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6551 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6552 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6553 cmirror_channel_0/VP outd_0/OutputN cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X6554 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6555 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6556 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6557 a_n17034_n701# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6558 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6559 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6560 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6561 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6562 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6563 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6564 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6565 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6566 cmirror_channel_0/VP outd_0/OutputP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X6567 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6568 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6569 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6570 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6571 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6572 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6573 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6574 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6575 isource_0/VM22D a_n35954_n3878# isource_0/VM3D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6576 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6577 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6578 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6579 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6580 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6581 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6582 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6583 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6584 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6585 outd_0/outd_stage1_0/isource_out outd_0/InputRef outd_0/V_da1_N outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6586 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6587 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6588 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6589 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6590 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6591 a_n17034_n701# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6592 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6593 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6594 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6595 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6596 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6597 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6598 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6599 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6600 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6601 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6602 cmirror_channel_0/TIA_I_Bias1 a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6603 tia_core_0/Out_2 outd_0/InputSignal tia_core_0/Input tia_core_0/Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6604 cmirror_channel_0/VP eigth_mirror_0/I_In a_n19500_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6605 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6606 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6607 tia_core_0/Input cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM5D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6608 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6609 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6610 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6611 cmirror_channel_0/VN isource_0/VM2D isource_0/VM2D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6612 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6613 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6614 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6615 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6616 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6617 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6618 tia_core_0/VM6D cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6619 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6620 isource_0/VM2D isource_0/VM2D cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6621 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6622 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6623 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6624 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6625 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6626 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6627 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6628 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6629 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6630 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6631 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6632 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6633 cmirror_channel_0/VN cmirror_channel_0/I_in_channel a_n6352_n5100# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6634 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6635 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6636 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6637 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6638 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6639 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6640 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6641 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6642 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6643 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6644 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6645 isource_0/VM11D isource_0/VM9D isource_0/VM8D isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6646 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6647 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6648 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6649 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6650 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6651 cmirror_channel_0/VN isource_0/VM2D isource_0/VM2D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6652 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6653 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6654 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6655 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6656 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6657 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6658 outd_0/V_da1_P cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
X6659 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6660 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6661 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6662 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6663 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6664 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6665 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6666 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6667 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6668 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6669 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6670 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6671 a_n20850_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6672 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6673 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6674 outd_0/outd_stage1_0/isource_out outd_0/InputRef outd_0/V_da1_N outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6675 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6676 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6677 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6678 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6679 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6680 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6681 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6682 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6683 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6684 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6685 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6686 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6687 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6688 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6689 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6690 cmirror_channel_0/VP outd_0/OutputP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X6691 outd_0/InputRef tia_core_0/VM39D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6692 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6693 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6694 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6695 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6696 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6697 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6698 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6699 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6700 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6701 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6702 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6703 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6704 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6705 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6706 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6707 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6708 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6709 tia_core_0/Input outd_0/InputSignal tia_core_0/Out_2 tia_core_0/Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6710 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6711 a_n11400_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6712 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6713 cmirror_channel_0/TIA_I_Bias1 a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6714 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6715 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6716 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6717 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6718 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6719 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6720 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6721 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6722 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6723 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6724 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6725 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6726 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6727 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6728 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6729 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6730 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6731 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6732 cmirror_channel_0/VP eigth_mirror_0/I_In a_n15450_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6733 cmirror_channel_0/VP cmirror_channel_0/VN tia_core_0/Out_2 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6734 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6735 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6736 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6737 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6738 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6739 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6740 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6741 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6742 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6743 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6744 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6745 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6746 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6747 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6748 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6749 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6750 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6751 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6752 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6753 cmirror_channel_0/VP eigth_mirror_0/I_In a_n11400_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6754 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6755 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6756 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6757 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6758 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6759 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6760 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6761 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6762 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6763 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6764 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6765 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6766 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6767 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6768 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6769 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6770 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6771 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6772 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6773 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6774 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6775 outd_0/outd_stage1_0/isource_out outd_0/InputSignal outd_0/V_da1_P outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6776 cmirror_channel_0/VP eigth_mirror_0/I_In a_n12750_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6777 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6778 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6779 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6780 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6781 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6782 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6783 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6784 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6785 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6786 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6787 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6788 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6789 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6790 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6791 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6792 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6793 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6794 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6795 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6796 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6797 tia_core_0/VM36D cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6798 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6799 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6800 cmirror_channel_0/VN isource_0/VM2D isource_0/VM2D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6801 tia_core_0/Input outd_0/InputSignal tia_core_0/Out_2 tia_core_0/Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6802 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6803 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6804 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6805 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6806 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6807 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6808 cmirror_channel_0/VP eigth_mirror_0/I_In a_n14100_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6809 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6810 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6811 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6812 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6813 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6814 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6815 tia_core_0/VM5D cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6816 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6817 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6818 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6819 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6820 isource_0/VM9D isource_0/VM9D isource_0/VM2D isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6821 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6822 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6823 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6824 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6825 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6826 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6827 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6828 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6829 isource_0/VM2D isource_0/VM2D cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6830 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6831 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6832 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6833 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6834 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6835 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6836 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6837 cmirror_channel_0/TIA_I_Bias1 a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6838 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6839 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6840 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6841 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6842 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6843 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6844 a_n12750_n11957# eigth_mirror_0/I_In cmirror_channel_0/I_in_channel cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6845 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6846 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6847 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6848 isource_0/VM3D a_n35954_n3878# isource_0/VM22D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6849 cmirror_channel_0/VP tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6850 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6851 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6852 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6853 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6854 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6855 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6856 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6857 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6858 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6859 a_n16464_n6284# a_n16994_n3852# cmirror_channel_0/VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X6860 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6861 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6862 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6863 outd_0/OutputN cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X6864 isource_0/VM8D isource_0/VM9D isource_0/VM11D isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6865 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6866 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6867 a_n11400_n11957# eigth_mirror_0/I_In eigth_mirror_0/I_In cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6868 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6869 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6870 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6871 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6872 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6873 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6874 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6875 tia_core_0/VM6D cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6876 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6877 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6878 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6879 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6880 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6881 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6882 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6883 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6884 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6885 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6886 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6887 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6888 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6889 cmirror_channel_0/A_Out_I_Bias a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6890 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6891 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6892 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6893 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6894 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6895 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6896 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6897 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6898 isource_0/VM9D isource_0/VM9D isource_0/VM2D isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6899 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6900 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6901 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6902 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6903 isource_0/VM11D isource_0/VM9D isource_0/VM8D isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6904 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6905 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6906 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6907 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6908 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6909 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6910 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6911 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6912 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6913 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6914 outd_0/InputRef tia_core_0/VM39D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6915 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6916 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6917 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6918 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6919 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6920 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6921 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6922 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6923 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6924 a_n35954_n3878# isource_0/VM22D eigth_mirror_0/I_In cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6925 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6926 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6927 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6928 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6929 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6930 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6931 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6932 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6933 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6934 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6935 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X6936 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6937 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6938 outd_0/OutputP cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X6939 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6940 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6941 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6942 a_n20054_26# a_n19524_2458# cmirror_channel_0/VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X6943 outd_0/V_da1_N outd_0/InputRef outd_0/outd_stage1_0/isource_out outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6944 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6945 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6946 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6947 cmirror_channel_0/VN cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM36D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6948 outd_0/outd_stage1_0/isource_out outd_0/InputSignal outd_0/V_da1_P outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6949 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6950 cmirror_channel_0/TIA_I_Bias1 a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6951 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6952 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6953 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6954 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6955 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6956 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6957 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6958 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6959 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6960 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6961 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6962 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6963 a_n4672_n5100# cmirror_channel_0/I_in_channel cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6964 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6965 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6966 outd_0/InputSignal tia_core_0/Input cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6967 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6968 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6969 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6970 outd_0/InputRef tia_core_0/VM39D tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6971 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6972 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6973 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6974 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6975 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6976 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6977 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6978 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6979 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6980 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6981 outd_0/OutputN cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X6982 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6983 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6984 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6985 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6986 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6987 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6988 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6989 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6990 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6991 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6992 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6993 cmirror_channel_0/TIA_I_Bias2 cmirror_channel_0/I_in_channel a_n4672_n5100# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X6994 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6995 a_n17034_n701# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6996 a_n17034_n701# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6997 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6998 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6999 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7000 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7001 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7002 a_n6352_n5100# cmirror_channel_0/I_in_channel cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7003 cmirror_channel_0/TIA_I_Bias1 tia_core_0/Disable_TIA cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7004 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7005 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7006 cmirror_channel_0/A_Out_I_Bias a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7007 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7008 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7009 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7010 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7011 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7012 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7013 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7014 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7015 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7016 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7017 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7018 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7019 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7020 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7021 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7022 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7023 cmirror_channel_0/VP eigth_mirror_0/I_In a_n18150_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7024 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7025 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7026 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7027 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7028 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7029 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7030 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7031 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7032 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7033 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7034 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7035 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7036 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7037 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7038 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7039 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7040 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7041 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7042 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7043 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7044 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7045 cmirror_channel_0/VN cmirror_channel_0/VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7046 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7047 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7048 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7049 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7050 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7051 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7052 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7053 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7054 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7055 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7056 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7057 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7058 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7059 a_n22200_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7060 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7061 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7062 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7063 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7064 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7065 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7066 cmirror_channel_0/VP eigth_mirror_0/I_In a_n19500_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7067 isource_0/VM8D isource_0/VM9D isource_0/VM11D isource_0/VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7068 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7069 isource_0/VM12G isource_0/VM14D cmirror_channel_0/VP isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7070 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7071 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7072 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X7073 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7074 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7075 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7076 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7077 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7078 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7079 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7080 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7081 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7082 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7083 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7084 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7085 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7086 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7087 outd_0/InputSignal tia_core_0/Input cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7088 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7089 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7090 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7091 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7092 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7093 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7094 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7095 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7096 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7097 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7098 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7099 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7100 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7101 outd_0/InputSignal tia_core_0/Input cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7102 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7103 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7104 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7105 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7106 cmirror_channel_0/VP outd_0/V_da2_N cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X7107 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7108 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7109 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7110 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7111 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7112 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7113 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7114 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7115 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7116 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7117 outd_0/outd_stage1_0/isource_out outd_0/InputRef outd_0/V_da1_N outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7118 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7119 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7120 a_n5250_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7121 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7122 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7123 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7124 cmirror_channel_0/VP cmirror_channel_0/VN tia_core_0/VM31D cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7125 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7126 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7127 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7128 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7129 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7130 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7131 isource_0/VM3D a_n35954_n3878# isource_0/VM22D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X7132 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7133 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7134 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7135 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7136 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7137 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7138 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7139 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7140 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7141 cmirror_channel_0/VP eigth_mirror_0/I_In a_n14100_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7142 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7143 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7144 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7145 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7146 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7147 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7148 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7149 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7150 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7151 cmirror_channel_0/VP outd_0/OutputN cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X7152 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7153 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7154 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7155 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7156 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7157 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7158 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7159 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7160 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7161 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7162 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7163 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7164 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7165 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7166 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7167 outd_0/InputRef tia_core_0/VM39D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7168 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7169 cmirror_channel_0/VP eigth_mirror_0/I_In a_n12750_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7170 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7171 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7172 tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__cap_var_lvt pd=0u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X7173 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7174 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7175 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7176 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7177 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7178 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7179 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7180 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7181 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7182 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7183 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7184 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7185 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7186 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7187 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7188 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7189 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7190 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7191 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7192 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7193 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7194 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7195 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7196 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7197 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7198 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7199 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7200 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7201 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7202 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7203 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7204 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7205 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7206 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7207 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7208 cmirror_channel_0/VN a_n18464_2458# cmirror_channel_0/VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X7209 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7210 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7211 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7212 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7213 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7214 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7215 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7216 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7217 outd_0/InputSignal tia_core_0/Input cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7218 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7219 isource_0/VM3D a_n35954_n3878# isource_0/VM22D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X7220 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7221 a_17268_7820# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7222 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7223 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7224 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7225 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7226 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7227 cmirror_channel_0/VP outd_0/OutputP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X7228 cmirror_channel_0/TIA_I_Bias1 cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM6D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7229 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7230 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7231 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7232 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7233 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7234 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7235 isource_0/VM2D isource_0/VM9D isource_0/VM9D isource_0/VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7236 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7237 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7238 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7239 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7240 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7241 tia_core_0/VM39D outd_0/InputRef tia_core_0/VM31D tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7242 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7243 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7244 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7245 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7246 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7247 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7248 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7249 tia_core_0/VM36D cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM39D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7250 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7251 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7252 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7253 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7254 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7255 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7256 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7257 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7258 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7259 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7260 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7261 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7262 cmirror_channel_0/VP isource_0/VM14D isource_0/VM12G isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7263 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7264 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7265 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7266 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7267 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7268 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7269 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7270 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7271 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7272 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7273 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7274 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7275 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7276 cmirror_channel_0/VN cmirror_channel_0/I_in_channel sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7277 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7278 isource_0/VM3G a_n21644_2458# cmirror_channel_0/VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X7279 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7280 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7281 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7282 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7283 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7284 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7285 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7286 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7287 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7288 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7289 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7290 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7291 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7292 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7293 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7294 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X7295 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7296 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7297 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7298 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7299 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7300 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7301 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7302 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7303 tia_core_0/VM31D outd_0/InputRef tia_core_0/VM39D tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7304 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7305 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7306 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7307 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7308 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7309 a_n22200_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7310 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7311 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7312 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7313 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7314 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7315 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7316 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7317 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7318 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7319 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7320 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7321 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7322 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7323 a_n17034_n2971# isource_0/VM8D cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7324 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7325 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7326 cmirror_channel_0/VN cmirror_channel_0/I_in_channel a_n6352_n5100# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7327 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7328 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7329 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7330 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7331 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7332 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7333 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7334 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7335 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7336 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7337 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7338 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7339 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7340 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7341 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7342 outd_0/outd_stage1_0/isource_out outd_0/InputSignal outd_0/V_da1_P outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7343 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7344 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7345 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7346 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7347 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7348 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7349 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7350 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7351 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7352 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7353 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7354 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7355 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7356 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7357 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7358 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7359 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7360 a_n17034_8339# isource_0/VM8D isource_0/VM9D cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X7361 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7362 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7363 outd_0/outd_stage1_0/isource_out cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7364 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7365 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7366 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7367 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7368 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7369 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7370 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7371 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7372 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7373 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7374 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7375 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7376 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7377 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7378 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7379 tia_core_0/VM31D cmirror_channel_0/VN cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7380 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7381 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7382 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7383 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7384 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7385 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7386 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7387 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7388 eigth_mirror_0/I_out_5 eigth_mirror_0/I_In a_n19500_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7389 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7390 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7391 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7392 a_n18150_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7393 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7394 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7395 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7396 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7397 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7398 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7399 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7400 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7401 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7402 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7403 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7404 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7405 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7406 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7407 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7408 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7409 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7410 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7411 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7412 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7413 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7414 cmirror_channel_0/VP isource_0/VM14D isource_0/VM12G isource_0/VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7415 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7416 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7417 isource_0/VM22D a_n35954_n3878# isource_0/VM3D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X7418 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7419 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7420 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7421 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7422 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7423 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7424 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7425 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7426 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7427 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7428 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7429 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7430 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7431 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7432 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7433 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7434 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7435 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7436 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7437 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17268_7820# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7438 outd_0/V_da1_N outd_0/InputRef outd_0/outd_stage1_0/isource_out outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7439 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7440 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7441 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7442 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7443 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7444 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7445 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7446 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7447 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7448 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7449 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7450 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7451 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7452 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7453 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7454 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7455 a_17890_7826# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage1_0/isource_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7456 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7457 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7458 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7459 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7460 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7461 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7462 isource_0/VM2D isource_0/VM2D cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X7463 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7464 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7465 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7466 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7467 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7468 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7469 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7470 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7471 cmirror_channel_0/A_Out_I_Bias a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7472 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7473 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7474 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7475 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7476 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7477 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7478 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7479 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7480 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7481 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7482 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7483 cmirror_channel_0/VN cmirror_channel_0/VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7484 cmirror_channel_0/VN isource_0/VM2D isource_0/VM2D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X7485 a_17890_7826# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7486 a_n17034_n701# isource_0/VM8D isource_0/VM14D cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X7487 a_n17034_n701# isource_0/VM8D isource_0/VM14D cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X7488 cmirror_channel_0/VP a_n5450_n3434# a_n3600_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7489 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7490 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7491 outd_0/V_da1_N cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
X7492 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7493 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7494 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7495 isource_0/VM22D a_n35954_n3878# isource_0/VM3D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X7496 outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7497 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7498 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7499 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7500 a_n15450_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7501 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7502 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7503 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7504 tia_core_0/VM31D outd_0/InputRef tia_core_0/VM39D tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7505 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7506 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7507 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7508 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7509 outd_0/V_da1_P cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
X7510 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7511 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7512 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7513 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7514 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7515 cmirror_channel_0/VP isource_0/VM8D a_n17034_8339# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7516 outd_0/V_da2_N outd_0/V_da1_N outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7517 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7518 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7519 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7520 a_n17034_n701# isource_0/VM8D isource_0/VM14D cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X7521 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7522 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7523 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7524 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7525 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7526 outd_0/OutputN cmirror_channel_0/VP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X7527 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7528 a_n22200_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7529 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7530 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7531 a_n14100_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7532 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7533 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7534 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7535 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7536 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7537 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7538 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7539 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7540 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7541 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7542 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7543 outd_0/InputSignal tia_core_0/Input cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7544 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7545 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7546 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7547 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM40D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7548 eigth_mirror_0/I_In isource_0/VM22D a_n35954_n3878# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7549 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7550 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7551 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7552 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7553 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7554 cmirror_channel_0/VP tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7555 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7556 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7557 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7558 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7559 outd_0/InputSignal tia_core_0/Input tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7560 outd_0/V_da1_P outd_0/InputSignal outd_0/outd_stage1_0/isource_out outd_0/outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7561 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7562 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7563 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7564 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7565 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7566 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7567 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7568 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7569 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7570 isource_0/VM11D isource_0/VM2D isource_0/VM12D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X7571 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7572 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7573 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7574 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7575 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7576 cmirror_channel_0/VP a_n5450_n3434# a_n5250_n3337# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7577 tia_core_0/VM31D outd_0/InputRef tia_core_0/VM39D tia_core_0/VM39D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7578 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7579 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7580 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7581 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7582 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7583 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7584 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7585 a_23060_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7586 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7587 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7588 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7589 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7590 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7591 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7592 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7593 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7594 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7595 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7596 cmirror_channel_0/VP eigth_mirror_0/I_In a_n14100_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7597 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7598 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7599 a_n17034_n701# isource_0/VM8D isource_0/VM14D cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X7600 isource_0/VM12D isource_0/VM2D isource_0/VM11D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X7601 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7602 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7603 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7604 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7605 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7606 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7607 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7608 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7609 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7610 outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7611 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7612 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7613 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7614 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7615 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7616 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7617 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7618 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7619 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7620 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7621 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7622 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7623 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_N outd_0/V_da2_N outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7624 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_P outd_0/OutputP outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7625 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7626 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7627 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7628 cmirror_channel_0/VP outd_0/OutputP cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X7629 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7630 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7631 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7632 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7633 cmirror_channel_0/VP eigth_mirror_0/I_In a_n12750_n11957# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7634 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7635 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7636 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7637 a_n18150_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7638 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7639 tia_core_0/VM40D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7640 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7641 a_n3600_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7642 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7643 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7644 isource_0/VM2D isource_0/VM2D cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X7645 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7646 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7647 cmirror_channel_0/VP a_n5450_n3434# a_n3320_n6897# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7648 tia_core_0/VM28D tia_core_0/Disable_TIA_B cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7649 outd_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7650 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7651 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7652 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7653 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_23060_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7654 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7655 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7656 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7657 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7658 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7659 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7660 outd_0/InputSignal tia_core_0/Input cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7661 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7662 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7663 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7664 cmirror_channel_0/VP isource_0/VM8D a_n17034_n701# cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7665 cmirror_channel_0/VN tia_core_0/Disable_TIA_B tia_core_0/VM28D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7666 tia_core_0/VM28D tia_core_0/Input outd_0/InputSignal cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7667 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7668 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7669 tia_core_0/VM36D cmirror_channel_0/TIA_I_Bias1 tia_core_0/VM39D cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7670 a_n16800_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7671 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7672 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7673 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7674 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7675 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7676 tia_core_0/VM40D tia_core_0/VM39D outd_0/InputRef cmirror_channel_0/VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7677 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7678 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7679 cmirror_channel_0/VP outd_0/OutputN cmirror_channel_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X7680 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7681 a_23060_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7682 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_17890_7826# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7683 tia_core_0/Out_2 outd_0/InputSignal tia_core_0/Input tia_core_0/Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X7684 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7685 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7686 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7687 a_n12750_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7688 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7689 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7690 outd_0/OutputN outd_0/V_da2_N outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7691 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7692 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7693 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7694 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7695 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7696 cmirror_channel_0/VN cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7697 a_37380_7026# cmirror_channel_0/A_Out_I_Bias outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7698 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out cmirror_channel_0/A_Out_I_Bias a_37380_7026# cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7699 outd_0/V_da2_P outd_0/V_da1_P outd_0/outd_stage2_0/cmirror_out outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7700 a_n5250_n3337# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7701 outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/V_da2_N outd_0/OutputN outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7702 a_n20850_n11957# eigth_mirror_0/I_In cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7703 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7704 a_n3320_n6897# a_n5450_n3434# cmirror_channel_0/VP cmirror_channel_0/VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7705 outd_0/outd_stage2_0/cmirror_out outd_0/V_da1_P outd_0/V_da2_P outd_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7706 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7707 outd_0/OutputP outd_0/V_da2_P outd_0/outd_stage3_0/outd_stage2_0/cmirror_out outd_0/outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7708 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7709 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7710 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7711 a_37380_7026# cmirror_channel_0/A_Out_I_Bias cmirror_channel_0/VN cmirror_channel_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
