magic
timestamp 1645191714
<< checkpaint >>
rect 0 -18910 8914 -260
<< pwell >>
rect 920 -17616 982 -17610
rect 920 -17610 922 -17540
rect 958 -14948 1020 -14942
rect 958 -14942 960 -14872
<< metal1 >>
rect 920 -18910 8519 -18876
rect 942 -18548 1042 -18348
rect 2652 -18548 2752 -18348
rect 4372 -18548 4472 -18348
rect 6092 -18548 6192 -18348
rect 7812 -18548 7912 -18348
rect 82 -18228 92 -18028
rect 172 -18228 182 -18028
rect 1802 -18228 1812 -18028
rect 1892 -18228 1902 -18028
rect 3512 -18228 3522 -18028
rect 3602 -18228 3612 -18028
rect 5232 -18228 5242 -18028
rect 5322 -18228 5332 -18028
rect 6942 -18228 6952 -18028
rect 7032 -18228 7042 -18028
rect 8662 -18228 8672 -18028
rect 8752 -18228 8762 -18028
rect 938 -17600 8425 -17566
rect 1032 -17566 8425 -17565
rect 958 -16242 8557 -16208
rect 980 -15880 1080 -15680
rect 2690 -15880 2790 -15680
rect 4410 -15880 4510 -15680
rect 6130 -15880 6230 -15680
rect 7850 -15880 7950 -15680
rect 120 -15560 130 -15360
rect 210 -15560 220 -15360
rect 1840 -15560 1850 -15360
rect 1930 -15560 1940 -15360
rect 3550 -15560 3560 -15360
rect 3640 -15560 3650 -15360
rect 5270 -15560 5280 -15360
rect 5360 -15560 5370 -15360
rect 6980 -15560 6990 -15360
rect 7070 -15560 7080 -15360
rect 8700 -15560 8710 -15360
rect 8790 -15560 8800 -15360
rect 976 -14932 8463 -14898
rect 1070 -14898 8463 -14897
<< via1 >>
rect 92 -18228 172 -18028
rect 1812 -18228 1892 -18028
rect 3522 -18228 3602 -18028
rect 5242 -18228 5322 -18028
rect 6952 -18228 7032 -18028
rect 8672 -18228 8752 -18028
rect 130 -15560 210 -15360
rect 1850 -15560 1930 -15360
rect 3560 -15560 3640 -15360
rect 5280 -15560 5360 -15360
rect 6990 -15560 7070 -15360
rect 8710 -15560 8790 -15360
<< metal2 >>
rect 952 -18558 1032 -18548
rect 2662 -18558 2742 -18548
rect 4382 -18558 4462 -18548
rect 6102 -18558 6182 -18548
rect 7822 -18558 7902 -18548
rect 952 -18348 1032 -18338
rect 2662 -18348 2742 -18338
rect 4382 -18348 4462 -18338
rect 6102 -18348 6182 -18338
rect 7822 -18348 7902 -18338
rect 92 -18238 172 -18228
rect 1812 -18238 1892 -18228
rect 3522 -18238 3602 -18228
rect 5242 -18238 5322 -18228
rect 6952 -18238 7032 -18228
rect 8672 -18238 8752 -18228
rect 172 -18228 1812 -18028
rect 1892 -18228 3522 -18028
rect 3602 -18228 5242 -18028
rect 5322 -18228 6952 -18028
rect 7032 -18228 8672 -18028
rect 8752 -18228 8762 -18028
rect 92 -18028 172 -18018
rect 1812 -18028 1892 -18018
rect 3522 -18028 3602 -18018
rect 5242 -18028 5322 -18018
rect 6952 -18028 7032 -18018
rect 8672 -18028 8752 -18018
rect 990 -15890 1070 -15880
rect 2700 -15890 2780 -15880
rect 4420 -15890 4500 -15880
rect 6140 -15890 6220 -15880
rect 7860 -15890 7940 -15880
rect 990 -15680 1070 -15670
rect 2700 -15680 2780 -15670
rect 4420 -15680 4500 -15670
rect 6140 -15680 6220 -15670
rect 7860 -15680 7940 -15670
rect 130 -15570 210 -15560
rect 1850 -15570 1930 -15560
rect 3560 -15570 3640 -15560
rect 5280 -15570 5360 -15560
rect 6990 -15570 7070 -15560
rect 8710 -15570 8790 -15560
rect 210 -15560 1850 -15360
rect 1930 -15560 3560 -15360
rect 3640 -15560 5280 -15360
rect 5360 -15560 6990 -15360
rect 7070 -15560 8710 -15360
rect 8790 -15560 8800 -15360
rect 130 -15360 210 -15350
rect 1850 -15360 1930 -15350
rect 3560 -15360 3640 -15350
rect 5280 -15360 5360 -15350
rect 6990 -15360 7070 -15350
rect 8710 -15360 8790 -15350
<< rmetal2 >>
rect 1032 -18548 2662 -18348
rect 2742 -18548 4382 -18348
rect 4462 -18548 6102 -18348
rect 6182 -18548 7822 -18348
rect 7902 -18548 8842 -18348
rect 1070 -15880 2700 -15680
rect 2780 -15880 4420 -15680
rect 4500 -15880 6140 -15680
rect 6220 -15880 7860 -15680
rect 7940 -15880 8880 -15680
use sky130_fd_pr__nfet_01v8_HH9N49 sky130_fd_pr__nfet_01v8_HH9N49_1
timestamp 1645191714
transform 1 0 4457 0 1 -2680
box -4457 -810 4457 810
use sky130_fd_pr__nfet_01v8_HH9N49 sky130_fd_pr__nfet_01v8_HH9N49_2
timestamp 1645191714
transform 1 0 4457 0 1 -1070
box -4457 -810 4457 810
use sky130_fd_pr__nfet_01v8_HH9N49 sky130_fd_pr__nfet_01v8_HH9N49_3
timestamp 1645191714
transform 1 0 4457 0 1 -4290
box -4457 -810 4457 810
use sky130_fd_pr__nfet_01v8_HH9N49 sky130_fd_pr__nfet_01v8_HH9N49_4
timestamp 1645191714
transform 1 0 4457 0 1 -5900
box -4457 -810 4457 810
use sky130_fd_pr__nfet_01v8_HH9N49 sky130_fd_pr__nfet_01v8_HH9N49_5
timestamp 1645191714
transform 1 0 4457 0 1 -7510
box -4457 -810 4457 810
use sky130_fd_pr__nfet_01v8_HH9N49 sky130_fd_pr__nfet_01v8_HH9N49_6
timestamp 1645191714
transform 1 0 4457 0 1 -9120
box -4457 -810 4457 810
use sky130_fd_pr__nfet_01v8_HH9N49 sky130_fd_pr__nfet_01v8_HH9N49_7
timestamp 1645191714
transform 1 0 4457 0 1 -10730
box -4457 -810 4457 810
use sky130_fd_pr__nfet_01v8_HH9N49 sky130_fd_pr__nfet_01v8_HH9N49_8
timestamp 1645191714
transform 1 0 4457 0 1 -12340
box -4457 -810 4457 810
use sky130_fd_pr__nfet_01v8_HH9N49 sky130_fd_pr__nfet_01v8_HH9N49_9
timestamp 1645191714
transform 1 0 4457 0 1 -13950
box -4457 -810 4457 810
use sky130_fd_pr__nfet_01v8_HH9N49 sky130_fd_pr__nfet_01v8_HH9N49_10
timestamp 1645191714
transform 1 0 4457 0 1 -15570
box -4457 -810 4457 810
<< end >>
