magic
tech sky130A
magscale 1 2
timestamp 1645802395
<< pwell >>
rect 122 552 1244 618
rect 122 42 1244 108
rect 130 -260 1640 -180
<< poly >>
rect 122 602 1244 618
rect 122 568 138 602
rect 172 568 330 602
rect 364 568 522 602
rect 556 568 714 602
rect 748 568 906 602
rect 940 568 1098 602
rect 1132 568 1244 602
rect 122 552 1244 568
rect 122 92 1244 108
rect 122 58 234 92
rect 268 58 426 92
rect 460 58 618 92
rect 652 58 810 92
rect 844 58 1002 92
rect 1036 58 1194 92
rect 1228 58 1244 92
rect 122 42 1244 58
<< polycont >>
rect 138 568 172 602
rect 330 568 364 602
rect 522 568 556 602
rect 714 568 748 602
rect 906 568 940 602
rect 1098 568 1132 602
rect 234 58 268 92
rect 426 58 460 92
rect 618 58 652 92
rect 810 58 844 92
rect 1002 58 1036 92
rect 1194 58 1228 92
<< locali >>
rect 122 568 138 602
rect 172 568 330 602
rect 364 568 522 602
rect 556 568 714 602
rect 748 568 906 602
rect 940 568 1098 602
rect 1132 568 1244 602
rect 122 58 234 92
rect 268 58 426 92
rect 460 58 618 92
rect 652 58 810 92
rect 844 58 1002 92
rect 1036 58 1194 92
rect 1228 58 1244 92
rect -20 -140 1390 -20
<< viali >>
rect 138 568 172 602
rect 330 568 364 602
rect 522 568 556 602
rect 714 568 748 602
rect 906 568 940 602
rect 1098 568 1132 602
rect 234 58 268 92
rect 426 58 460 92
rect 618 58 652 92
rect 810 58 844 92
rect 1002 58 1036 92
rect 1194 58 1228 92
<< metal1 >>
rect 120 602 1440 630
rect 120 568 138 602
rect 172 568 330 602
rect 364 568 522 602
rect 556 568 714 602
rect 748 568 906 602
rect 940 568 1098 602
rect 1132 568 1440 602
rect 120 560 1440 568
rect 167 370 177 530
rect 229 370 239 530
rect 359 370 369 530
rect 421 370 431 530
rect 551 370 561 530
rect 613 370 623 530
rect 743 370 753 530
rect 805 370 815 530
rect 935 370 945 530
rect 997 370 1007 530
rect 1127 370 1137 530
rect 1189 370 1199 530
rect 71 130 81 290
rect 133 130 143 290
rect 263 130 273 290
rect 325 130 335 290
rect 455 130 465 290
rect 517 130 527 290
rect 647 130 657 290
rect 709 130 719 290
rect 839 130 849 290
rect 901 130 911 290
rect 1031 130 1041 290
rect 1093 130 1103 290
rect 1223 130 1233 290
rect 1285 130 1295 290
rect 1330 100 1440 560
rect 120 92 1440 100
rect 120 58 234 92
rect 268 58 426 92
rect 460 58 618 92
rect 652 58 810 92
rect 844 58 1002 92
rect 1036 58 1194 92
rect 1228 58 1440 92
rect 120 30 1440 58
rect 1310 -180 1440 30
rect 130 -260 1640 -180
rect 329 -450 339 -290
rect 391 -450 401 -290
rect 845 -450 855 -290
rect 907 -450 917 -290
rect 1361 -450 1371 -290
rect 1423 -450 1430 -290
rect 71 -690 81 -530
rect 133 -690 143 -530
rect 587 -690 597 -530
rect 649 -690 659 -530
rect 1103 -690 1113 -530
rect 1165 -690 1175 -530
rect 1480 -720 1570 -260
rect 1619 -690 1629 -530
rect 1681 -690 1691 -530
rect 70 -800 1690 -720
<< via1 >>
rect 177 370 229 530
rect 369 370 421 530
rect 561 370 613 530
rect 753 370 805 530
rect 945 370 997 530
rect 1137 370 1189 530
rect 81 130 133 290
rect 273 130 325 290
rect 465 130 517 290
rect 657 130 709 290
rect 849 130 901 290
rect 1041 130 1093 290
rect 1233 130 1285 290
rect 339 -450 391 -290
rect 855 -450 907 -290
rect 1371 -450 1423 -290
rect 81 -690 133 -530
rect 597 -690 649 -530
rect 1113 -690 1165 -530
rect 1629 -690 1681 -530
<< metal2 >>
rect 170 530 1200 540
rect 170 370 177 530
rect 229 370 369 530
rect 421 370 561 530
rect 613 370 753 530
rect 805 370 945 530
rect 997 370 1137 530
rect 1189 370 1200 530
rect 170 360 1200 370
rect 80 290 1430 300
rect 80 130 81 290
rect 133 130 273 290
rect 325 130 465 290
rect 517 130 657 290
rect 709 130 849 290
rect 901 130 1041 290
rect 1093 130 1233 290
rect 1285 130 1430 290
rect 80 120 1430 130
rect 1130 -260 1430 120
rect 320 -290 1430 -260
rect 320 -450 339 -290
rect 391 -450 855 -290
rect 907 -450 1371 -290
rect 1423 -450 1430 -290
rect 320 -460 1430 -450
rect 70 -530 1690 -520
rect 70 -690 81 -530
rect 133 -690 597 -530
rect 649 -690 1113 -530
rect 1165 -690 1629 -530
rect 1681 -690 1690 -530
rect 70 -700 1690 -690
use sky130_fd_pr__nfet_01v8_854667  sky130_fd_pr__nfet_01v8_854667_0
timestamp 1645802395
transform 1 0 881 0 1 -490
box -941 -410 941 410
use sky130_fd_pr__nfet_01v8_F8VELN  sky130_fd_pr__nfet_01v8_F8VELN_0
timestamp 1645801865
transform 1 0 683 0 1 330
box -743 -410 743 410
<< end >>
