magic
tech sky130A
magscale 1 2
timestamp 1646921651
<< nwell >>
rect -9230 1690 -1970 1730
rect -8600 1110 -8450 1690
rect -7870 1110 -7720 1690
rect -7130 1110 -6980 1690
rect -6400 1110 -6250 1690
rect -5670 1110 -5520 1690
rect -4940 1110 -4790 1690
rect -4210 1110 -4060 1690
rect -3470 1080 -3330 1690
rect -2740 1060 -2600 1690
rect -2010 1080 -1970 1690
<< pwell >>
rect -9370 1830 -1830 1870
rect -8600 300 -8440 930
rect -7870 300 -7710 930
rect -7140 300 -6980 930
rect -6400 290 -6240 920
rect -5670 300 -5510 930
rect -4940 290 -4780 920
rect -4210 290 -4050 920
rect -3480 280 -3320 910
<< locali >>
rect -9370 1830 -1830 1870
rect -9370 980 -9320 1830
rect -9230 1720 -1970 1730
rect -9230 1070 -9220 1720
rect -1980 1070 -1970 1720
rect -9230 1060 -1970 1070
rect -9370 270 -9340 980
rect -1880 970 -1830 1830
rect -1870 270 -1830 970
rect -9370 260 -1830 270
<< viali >>
rect -9220 1660 -1980 1720
rect -9220 1130 -9170 1660
rect -8620 1130 -8440 1660
rect -7890 1130 -7710 1660
rect -7150 1130 -6970 1660
rect -6420 1130 -6240 1660
rect -5690 1130 -5510 1660
rect -4960 1130 -4780 1660
rect -4220 1130 -4040 1660
rect -3490 1130 -3310 1660
rect -2760 1130 -2580 1660
rect -2030 1130 -1980 1660
rect -9220 1070 -1980 1130
rect -9340 970 -9170 980
rect -8610 970 -8440 980
rect -7880 970 -7710 980
rect -7150 970 -6980 980
rect -6410 970 -6240 980
rect -5680 970 -5510 980
rect -4950 970 -4780 980
rect -4220 970 -4050 980
rect -3490 970 -3320 980
rect -2760 970 -2590 980
rect -9340 870 -1870 970
rect -9340 330 -9170 870
rect -8610 330 -8440 870
rect -7880 330 -7710 870
rect -7150 330 -6980 870
rect -6410 330 -6240 870
rect -5680 330 -5510 870
rect -4950 330 -4780 870
rect -4220 330 -4050 870
rect -3490 330 -3320 870
rect -2760 330 -2590 870
rect -2020 330 -1870 870
rect -9340 270 -1870 330
<< metal1 >>
rect -9290 1720 -1910 1990
rect -9290 1070 -9220 1720
rect -9170 1654 -8620 1660
rect -9170 1136 -9160 1654
rect -9090 1210 -9080 1590
rect -8700 1210 -8690 1590
rect -8630 1136 -8620 1654
rect -9170 1130 -8620 1136
rect -8440 1654 -7890 1660
rect -8440 1136 -8430 1654
rect -8360 1210 -8350 1586
rect -7974 1210 -7964 1586
rect -7900 1136 -7890 1654
rect -8440 1130 -7890 1136
rect -7710 1654 -7150 1660
rect -7710 1136 -7700 1654
rect -7630 1200 -7620 1576
rect -7244 1200 -7234 1576
rect -7160 1136 -7150 1654
rect -7710 1130 -7150 1136
rect -6970 1654 -6420 1660
rect -6970 1136 -6960 1654
rect -6900 1200 -6890 1576
rect -6514 1200 -6504 1576
rect -6430 1136 -6420 1654
rect -6970 1130 -6420 1136
rect -6240 1654 -5690 1660
rect -6240 1136 -6230 1654
rect -6170 1200 -6160 1576
rect -5784 1200 -5774 1576
rect -5700 1136 -5690 1654
rect -6240 1130 -5690 1136
rect -5510 1654 -4960 1660
rect -5510 1136 -5500 1654
rect -5440 1200 -5430 1576
rect -5054 1200 -5044 1576
rect -4970 1136 -4960 1654
rect -5510 1130 -4960 1136
rect -4780 1654 -4220 1660
rect -4780 1136 -4770 1654
rect -4700 1210 -4690 1586
rect -4314 1210 -4304 1586
rect -4230 1136 -4220 1654
rect -4780 1130 -4220 1136
rect -4040 1654 -3490 1660
rect -4040 1136 -4030 1654
rect -3970 1210 -3960 1586
rect -3584 1210 -3574 1586
rect -3500 1136 -3490 1654
rect -4040 1130 -3490 1136
rect -3310 1654 -2760 1660
rect -3310 1136 -3300 1654
rect -3230 1210 -3220 1586
rect -2844 1210 -2834 1586
rect -2770 1136 -2760 1654
rect -3310 1130 -2760 1136
rect -2580 1654 -2030 1660
rect -2580 1136 -2570 1654
rect -2500 1210 -2490 1586
rect -2114 1210 -2104 1586
rect -2040 1136 -2030 1654
rect -2580 1130 -2030 1136
rect -1980 1070 -1910 1720
rect -9290 1064 -1910 1070
rect -9290 1060 -9160 1064
rect -8630 1060 -8430 1064
rect -7900 1060 -7700 1064
rect -7160 1060 -6960 1064
rect -6430 1060 -6230 1064
rect -5700 1060 -5500 1064
rect -4970 1060 -4770 1064
rect -4230 1060 -4030 1064
rect -3500 1060 -3300 1064
rect -2770 1060 -2570 1064
rect -2040 1060 -1910 1064
rect -9226 1058 -9164 1060
rect -8626 1058 -8434 1060
rect -7896 1058 -7704 1060
rect -7156 1058 -6964 1060
rect -6426 1058 -6234 1060
rect -5696 1058 -5504 1060
rect -4966 1058 -4774 1060
rect -4226 1058 -4034 1060
rect -3496 1058 -3304 1060
rect -2766 1058 -2574 1060
rect -2036 1058 -1974 1060
rect -9346 990 -9164 992
rect -8616 990 -8434 992
rect -7886 990 -7704 992
rect -7156 990 -6974 992
rect -6416 990 -6234 992
rect -5686 990 -5504 992
rect -4956 990 -4774 992
rect -4226 990 -4044 992
rect -3496 990 -3314 992
rect -2766 990 -2584 992
rect -9350 980 -9160 990
rect -9350 976 -9340 980
rect -9352 864 -9340 976
rect -9170 976 -9160 980
rect -8620 980 -8430 990
rect -8620 976 -8610 980
rect -9170 970 -8610 976
rect -8440 976 -8430 980
rect -7890 980 -7700 990
rect -7890 976 -7880 980
rect -8440 970 -7880 976
rect -7710 976 -7700 980
rect -7160 980 -6970 990
rect -7160 976 -7150 980
rect -7710 970 -7150 976
rect -6980 976 -6970 980
rect -6420 980 -6230 990
rect -6420 976 -6410 980
rect -6980 970 -6410 976
rect -6240 976 -6230 980
rect -5690 980 -5500 990
rect -5690 976 -5680 980
rect -6240 970 -5680 976
rect -5510 976 -5500 980
rect -4960 980 -4770 990
rect -4960 976 -4950 980
rect -5510 970 -4950 976
rect -4780 976 -4770 980
rect -4230 980 -4030 990
rect -4230 976 -4220 980
rect -4780 970 -4220 976
rect -4050 976 -4030 980
rect -3500 980 -3300 990
rect -3500 976 -3490 980
rect -4050 970 -3490 976
rect -3320 976 -3300 980
rect -2770 980 -2570 990
rect -2026 980 -1864 982
rect -2770 976 -2760 980
rect -3320 970 -2760 976
rect -2590 976 -2570 980
rect -2030 976 -1860 980
rect -2590 970 -1858 976
rect -9350 336 -9340 864
rect -9352 270 -9340 336
rect -9170 864 -8610 870
rect -9170 336 -9160 864
rect -9090 410 -9080 790
rect -8700 410 -8690 790
rect -8620 336 -8610 864
rect -9170 330 -8610 336
rect -8440 864 -7880 870
rect -8440 336 -8430 864
rect -8360 410 -8350 790
rect -7970 410 -7960 790
rect -7890 336 -7880 864
rect -8440 330 -7880 336
rect -7710 864 -7150 870
rect -7710 336 -7700 864
rect -7630 410 -7620 790
rect -7240 410 -7230 790
rect -7160 336 -7150 864
rect -7710 330 -7150 336
rect -6980 864 -6410 870
rect -6980 336 -6970 864
rect -6900 410 -6890 790
rect -6510 410 -6500 790
rect -6420 336 -6410 864
rect -6980 330 -6410 336
rect -6240 864 -5680 870
rect -6240 336 -6230 864
rect -6170 410 -6160 790
rect -5780 410 -5770 790
rect -5690 336 -5680 864
rect -6240 330 -5680 336
rect -5510 864 -4950 870
rect -5510 336 -5500 864
rect -5430 410 -5420 790
rect -5040 410 -5030 790
rect -4960 336 -4950 864
rect -5510 330 -4950 336
rect -4780 864 -4220 870
rect -4780 336 -4770 864
rect -4700 410 -4690 790
rect -4310 410 -4300 790
rect -4230 336 -4220 864
rect -4780 330 -4220 336
rect -4050 864 -3490 870
rect -4050 336 -4030 864
rect -3970 410 -3960 790
rect -3580 410 -3570 790
rect -3500 336 -3490 864
rect -4050 330 -3490 336
rect -3320 864 -2760 870
rect -3320 336 -3300 864
rect -3240 410 -3230 790
rect -2850 410 -2840 790
rect -2770 336 -2760 864
rect -3320 330 -2760 336
rect -2590 864 -2020 870
rect -2590 336 -2570 864
rect -2500 410 -2490 790
rect -2110 410 -2100 790
rect -2030 336 -2020 864
rect -2590 330 -2020 336
rect -1870 864 -1858 970
rect -1870 336 -1860 864
rect -1870 270 -1858 336
rect -9352 264 -1858 270
rect -9350 60 -1860 264
<< via1 >>
rect -9080 1210 -8700 1590
rect -8350 1210 -7974 1586
rect -7620 1200 -7244 1576
rect -6890 1200 -6514 1576
rect -6160 1200 -5784 1576
rect -5430 1200 -5054 1576
rect -4690 1210 -4314 1586
rect -3960 1210 -3584 1586
rect -3220 1210 -2844 1586
rect -2490 1210 -2114 1586
rect -9080 410 -8700 790
rect -8350 410 -7970 790
rect -7620 410 -7240 790
rect -6890 410 -6510 790
rect -6160 410 -5780 790
rect -5420 410 -5040 790
rect -4690 410 -4310 790
rect -3960 410 -3580 790
rect -3230 410 -2850 790
rect -2490 410 -2110 790
<< metal2 >>
rect -9090 1590 -2100 1600
rect -9090 1210 -9080 1590
rect -8700 1586 -2100 1590
rect -8700 1210 -8350 1586
rect -7974 1576 -4690 1586
rect -7974 1210 -7620 1576
rect -9090 1200 -7620 1210
rect -7244 1200 -6890 1576
rect -6514 1200 -6160 1576
rect -5784 1200 -5430 1576
rect -5054 1210 -4690 1576
rect -4314 1210 -3960 1586
rect -3584 1210 -3220 1586
rect -2844 1210 -2490 1586
rect -2114 1210 -2100 1586
rect -5054 1200 -2100 1210
rect -9090 790 -2100 1200
rect -9090 410 -9080 790
rect -8700 410 -8350 790
rect -7970 410 -7620 790
rect -7240 410 -6890 790
rect -6510 410 -6160 790
rect -5780 410 -5420 790
rect -5040 410 -4690 790
rect -4310 410 -3960 790
rect -3580 410 -3230 790
rect -2850 410 -2490 790
rect -2110 410 -2100 790
rect -9090 400 -2100 410
use sky130_fd_pr__diode_pd2nw_05v5_33C8ED  sky130_fd_pr__diode_pd2nw_05v5_33C8ED_0
timestamp 1646921651
transform 1 0 -5599 0 1 1395
box -3770 -476 3770 476
use sky130_fd_pr__diode_pw2nd_05v5_T9UBGD  sky130_fd_pr__diode_pw2nd_05v5_T9UBGD_0
timestamp 1646921651
transform 1 0 -5598 0 1 598
box -3632 -338 3632 338
<< end >>
