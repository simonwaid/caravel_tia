magic
tech sky130A
magscale 1 2
timestamp 1646921651
<< dnwell >>
rect 60 8030 12100 9910
<< nwell >>
rect -20 9704 12180 9990
rect -20 8236 266 9704
rect 11894 8236 12180 9704
rect -20 7950 12180 8236
<< pwell >>
rect 3000 11360 3030 11440
<< nsubdiff >>
rect 17 9933 12143 9953
rect 17 9899 97 9933
rect 12063 9899 12143 9933
rect 17 9879 12143 9899
rect 17 9873 91 9879
rect 17 8067 37 9873
rect 71 8067 91 9873
rect 17 8061 91 8067
rect 12069 9873 12143 9879
rect 12069 8067 12089 9873
rect 12123 8067 12143 9873
rect 12069 8061 12143 8067
rect 17 8041 12143 8061
rect 17 8007 97 8041
rect 12063 8007 12143 8041
rect 17 7987 12143 8007
<< nsubdiffcont >>
rect 97 9899 12063 9933
rect 37 8067 71 9873
rect 12089 8067 12123 9873
rect 97 8007 12063 8041
<< locali >>
rect 1640 12030 1740 13940
rect 3100 12030 3200 13940
rect 4570 12030 4670 13940
rect 6030 12030 6130 13940
rect 7490 12030 7600 13940
rect 8960 12030 9070 13940
rect 10430 12030 10540 13940
rect 11880 12030 12160 13940
rect 250 11940 12160 12030
rect 1640 10740 1740 11940
rect 1630 10700 1740 10740
rect 1630 10040 1730 10700
rect 3100 10040 3200 11940
rect 4570 10750 4670 11940
rect 4560 10040 4670 10750
rect 6030 10750 6130 11940
rect 6030 10040 6140 10750
rect 7490 10040 7600 11940
rect 8960 10040 9070 11940
rect 10430 10750 10540 11940
rect 10420 10700 10540 10750
rect 10420 10040 10530 10700
rect 11880 10300 12160 11940
rect 11880 10040 12510 10300
rect 50 9933 1460 9950
rect 1950 9933 4350 9950
rect 4900 9933 7270 9950
rect 7820 9933 10190 9950
rect 10740 9933 12120 9950
rect 37 9899 97 9933
rect 12063 9899 12123 9933
rect 37 9873 71 9899
rect 12089 9873 12123 9899
rect 300 9620 11860 9690
rect 300 8320 350 9620
rect 1630 9250 1730 9620
rect 1630 8320 1730 8690
rect 3020 8320 3280 9620
rect 4560 9250 4660 9620
rect 4560 8320 4660 8690
rect 5950 8320 6210 9620
rect 7490 9250 7590 9620
rect 7490 8320 7590 8690
rect 8880 8320 9140 9620
rect 10420 9250 10520 9620
rect 10420 8320 10520 8690
rect 11810 8320 11860 9620
rect 300 8250 11860 8320
rect 37 8041 71 8067
rect 12089 8041 12123 8067
rect 37 8007 97 8041
rect 12063 8007 12123 8041
rect 12250 7990 12510 10040
rect 12250 7900 13370 7990
rect 12420 7890 13370 7900
rect 13210 5200 13360 7890
<< viali >>
rect 1460 9933 1950 9970
rect 4350 9933 4900 9960
rect 7270 9933 7820 9960
rect 10190 9933 10740 9960
rect 1460 9899 1950 9933
rect 4350 9899 4900 9933
rect 7270 9899 7820 9933
rect 10190 9899 10740 9933
rect 1460 9880 1950 9899
rect 4350 9880 4900 9899
rect 7270 9880 7820 9899
rect 10190 9880 10740 9899
rect 1620 8690 1750 9250
rect 4550 8690 4680 9250
rect 7480 8690 7610 9250
rect 10410 8690 10540 9250
<< metal1 >>
rect 1100 13380 1110 13820
rect 2260 13380 2270 13820
rect 4030 13380 4040 13820
rect 5190 13380 5200 13820
rect 6960 13380 6970 13820
rect 8120 13380 8130 13820
rect 9890 13380 9900 13820
rect 11050 13380 11060 13820
rect 370 11400 380 12580
rect 1010 11400 1020 12580
rect 2350 11400 2360 12580
rect 2990 11400 3000 12580
rect 3300 11400 3310 12580
rect 3940 11400 3950 12580
rect 5280 11400 5290 12580
rect 5920 11400 5930 12580
rect 6230 11400 6240 12580
rect 6870 11400 6880 12580
rect 8210 11400 8220 12580
rect 8850 11400 8860 12580
rect 9160 11400 9170 12580
rect 9800 11400 9810 12580
rect 11140 11400 11150 12580
rect 11780 11400 11790 12580
rect 1100 10160 1110 10600
rect 2260 10160 2270 10600
rect 4030 10160 4040 10600
rect 5190 10160 5200 10600
rect 6960 10160 6970 10600
rect 8120 10160 8130 10600
rect 9890 10160 9900 10600
rect 11050 10160 11060 10600
rect 1460 9976 1950 10160
rect 1448 9970 1962 9976
rect 1448 9880 1460 9970
rect 1950 9880 1962 9970
rect 4350 9966 4900 10160
rect 7270 9966 7820 10160
rect 10190 9966 10740 10160
rect 1448 9874 1962 9880
rect 4338 9960 4912 9966
rect 4338 9880 4350 9960
rect 4900 9880 4912 9960
rect 4338 9874 4912 9880
rect 7258 9960 7832 9966
rect 7258 9880 7270 9960
rect 7820 9880 7832 9960
rect 7258 9874 7832 9880
rect 10178 9960 10752 9966
rect 10178 9880 10190 9960
rect 10740 9880 10752 9960
rect 10178 9874 10752 9880
rect 330 9510 1510 9570
rect 1850 9510 3040 9570
rect 330 9050 400 9510
rect 1614 9250 1756 9262
rect 330 9040 1510 9050
rect 250 8900 260 9040
rect 390 8990 1510 9040
rect 390 8950 400 8990
rect 390 8900 1510 8950
rect 330 8890 1510 8900
rect 330 8430 400 8890
rect 1610 8690 1620 9250
rect 1750 8690 1760 9250
rect 2970 9040 3040 9510
rect 3260 9510 4440 9570
rect 4780 9510 5970 9570
rect 3260 9050 3330 9510
rect 4544 9250 4686 9262
rect 3260 9040 4440 9050
rect 1850 8980 2980 9040
rect 2970 8950 2980 8980
rect 1850 8900 2980 8950
rect 3110 8900 3120 9040
rect 3180 8900 3190 9040
rect 3320 8990 4440 9040
rect 3320 8950 3330 8990
rect 3320 8900 4440 8950
rect 1850 8890 3040 8900
rect 1614 8678 1756 8690
rect 2970 8430 3040 8890
rect 330 8370 1510 8430
rect 1850 8370 3040 8430
rect 3260 8890 4440 8900
rect 3260 8430 3330 8890
rect 4540 8690 4550 9250
rect 4680 8690 4690 9250
rect 5900 9040 5970 9510
rect 6190 9510 7370 9570
rect 7710 9510 8900 9570
rect 6190 9050 6260 9510
rect 7474 9250 7616 9262
rect 6190 9040 7370 9050
rect 4780 8980 5910 9040
rect 5900 8950 5910 8980
rect 4780 8900 5910 8950
rect 6040 8900 6050 9040
rect 6110 8900 6120 9040
rect 6250 8990 7370 9040
rect 6250 8950 6260 8990
rect 6250 8900 7370 8950
rect 4780 8890 5970 8900
rect 4544 8678 4686 8690
rect 5900 8430 5970 8890
rect 3260 8370 4440 8430
rect 4780 8370 5970 8430
rect 6190 8890 7370 8900
rect 6190 8430 6260 8890
rect 7470 8690 7480 9250
rect 7610 8690 7620 9250
rect 8830 9040 8900 9510
rect 9120 9510 10300 9570
rect 10640 9510 11830 9570
rect 9120 9050 9190 9510
rect 10404 9250 10546 9262
rect 9120 9040 10300 9050
rect 7710 8980 8840 9040
rect 8830 8950 8840 8980
rect 7710 8900 8840 8950
rect 8970 8900 8980 9040
rect 9040 8910 9050 9040
rect 9180 8990 10300 9040
rect 9180 8950 9190 8990
rect 9180 8910 10300 8950
rect 7710 8890 8900 8900
rect 7474 8678 7616 8690
rect 8830 8430 8900 8890
rect 6190 8370 7370 8430
rect 7710 8370 8900 8430
rect 9120 8890 10300 8910
rect 9120 8430 9190 8890
rect 10400 8690 10410 9250
rect 10540 8690 10550 9250
rect 11760 9040 11830 9510
rect 10640 8980 11770 9040
rect 11760 8950 11770 8980
rect 10640 8900 11770 8950
rect 11900 8900 11910 9040
rect 10640 8890 11830 8900
rect 10404 8678 10546 8690
rect 11760 8430 11830 8890
rect 9120 8370 10300 8430
rect 10640 8370 11830 8430
<< via1 >>
rect 1110 13380 2260 13820
rect 4040 13380 5190 13820
rect 6970 13380 8120 13820
rect 9900 13380 11050 13820
rect 380 11400 1010 12580
rect 2360 11400 2990 12580
rect 3310 11400 3940 12580
rect 5290 11400 5920 12580
rect 6240 11400 6870 12580
rect 8220 11400 8850 12580
rect 9170 11400 9800 12580
rect 11150 11400 11780 12580
rect 1110 10160 2260 10600
rect 4040 10160 5190 10600
rect 6970 10160 8120 10600
rect 9900 10160 11050 10600
rect 260 8900 390 9040
rect 1620 8690 1750 9250
rect 2980 8900 3110 9040
rect 3190 8900 3320 9040
rect 4550 8690 4680 9250
rect 5910 8900 6040 9040
rect 6120 8900 6250 9040
rect 7480 8690 7610 9250
rect 8840 8900 8970 9040
rect 9050 8910 9180 9040
rect 10410 8690 10540 9250
rect 11770 8900 11900 9040
<< metal2 >>
rect 1110 13820 2260 13830
rect 1110 13370 2260 13380
rect 4040 13820 5190 13830
rect 4040 13370 5190 13380
rect 6970 13820 8120 13830
rect 6970 13370 8120 13380
rect 9900 13820 11050 13830
rect 9900 13370 11050 13380
rect 380 12580 1010 12590
rect 380 11390 1010 11400
rect 2360 12580 2990 12590
rect 2360 11390 2990 11400
rect 3310 12580 3940 12590
rect 3310 11390 3940 11400
rect 5290 12580 5920 12590
rect 5290 11390 5920 11400
rect 6240 12580 6870 12590
rect 6240 11390 6870 11400
rect 8220 12580 8850 12590
rect 8220 11390 8850 11400
rect 9170 12580 9800 12590
rect 9170 11390 9800 11400
rect 11150 12580 11780 12590
rect 11150 11390 11780 11400
rect 1110 10600 2260 10610
rect 1110 10150 2260 10160
rect 4040 10600 5190 10610
rect 4040 10150 5190 10160
rect 6970 10600 8120 10610
rect 6970 10150 8120 10160
rect 9900 10600 11050 10610
rect 9900 10150 11050 10160
rect -20 9520 11910 9690
rect 250 9040 400 9520
rect 440 9470 1450 9480
rect 440 9330 450 9470
rect 1000 9330 1450 9470
rect 440 9320 1450 9330
rect 1910 9470 2930 9480
rect 1910 9330 2370 9470
rect 2920 9330 2930 9470
rect 1910 9320 2930 9330
rect 1620 9250 1750 9260
rect 540 9230 1620 9240
rect 1750 9230 2830 9240
rect 540 9090 1100 9230
rect 2270 9090 2830 9230
rect 540 9080 1620 9090
rect 250 8900 260 9040
rect 390 8900 400 9040
rect 250 8890 400 8900
rect 540 8850 1620 8860
rect 1750 9080 2830 9090
rect 2980 9040 3110 9050
rect 3180 9040 3330 9520
rect 3370 9470 4380 9480
rect 3370 9330 3380 9470
rect 3930 9330 4380 9470
rect 3370 9320 4380 9330
rect 4840 9470 5860 9480
rect 4840 9330 5300 9470
rect 5850 9330 5860 9470
rect 4840 9320 5860 9330
rect 4550 9250 4680 9260
rect 3470 9230 4550 9240
rect 4680 9230 5760 9240
rect 3470 9090 4030 9230
rect 5200 9090 5760 9230
rect 3470 9080 4550 9090
rect 2970 8900 2980 9040
rect 3110 8900 3120 9040
rect 1750 8850 2830 8860
rect 540 8710 1100 8850
rect 2270 8710 2830 8850
rect 540 8700 1620 8710
rect 1750 8700 2830 8710
rect 1620 8680 1750 8690
rect 440 8610 1450 8620
rect 440 8470 450 8610
rect 1000 8470 1450 8610
rect 440 8460 1450 8470
rect 1910 8610 2930 8620
rect 1910 8470 2370 8610
rect 2920 8470 2930 8610
rect 1910 8460 2930 8470
rect 2970 8420 3120 8900
rect 3180 8900 3190 9040
rect 3320 8900 3330 9040
rect 3180 8890 3330 8900
rect 3470 8850 4550 8860
rect 4680 9080 5760 9090
rect 5910 9040 6040 9050
rect 6110 9040 6260 9520
rect 6300 9470 7310 9480
rect 6300 9330 6310 9470
rect 6860 9330 7310 9470
rect 6300 9320 7310 9330
rect 7770 9470 8790 9480
rect 7770 9330 8230 9470
rect 8780 9330 8790 9470
rect 7770 9320 8790 9330
rect 7480 9250 7610 9260
rect 6400 9230 7480 9240
rect 7610 9230 8690 9240
rect 6400 9090 6960 9230
rect 8130 9090 8690 9230
rect 6400 9080 7480 9090
rect 5900 8900 5910 9040
rect 6040 8900 6050 9040
rect 4680 8850 5760 8860
rect 3470 8710 4030 8850
rect 5200 8710 5760 8850
rect 3470 8700 4550 8710
rect 4680 8700 5760 8710
rect 4550 8680 4680 8690
rect 3370 8610 4380 8620
rect 3370 8470 3380 8610
rect 3930 8470 4380 8610
rect 3370 8460 4380 8470
rect 4840 8610 5860 8620
rect 4840 8470 5300 8610
rect 5850 8470 5860 8610
rect 4840 8460 5860 8470
rect 5900 8420 6050 8900
rect 6110 8900 6120 9040
rect 6250 8900 6260 9040
rect 6110 8890 6260 8900
rect 6400 8850 7480 8860
rect 7610 9080 8690 9090
rect 8840 9040 8970 9050
rect 9040 9040 9190 9520
rect 9230 9470 10240 9480
rect 9230 9330 9240 9470
rect 9790 9330 10240 9470
rect 9230 9320 10240 9330
rect 10700 9470 11720 9480
rect 10700 9330 11160 9470
rect 11710 9330 11720 9470
rect 10700 9320 11720 9330
rect 10410 9250 10540 9260
rect 9330 9230 10410 9240
rect 10540 9230 11620 9240
rect 9330 9090 9890 9230
rect 11060 9090 11620 9230
rect 9330 9080 10410 9090
rect 8830 8900 8840 9040
rect 8970 8900 8980 9040
rect 9040 8910 9050 9040
rect 9180 8910 9190 9040
rect 9040 8900 9190 8910
rect 7610 8850 8690 8860
rect 6400 8710 6960 8850
rect 8130 8710 8690 8850
rect 6400 8700 7480 8710
rect 7610 8700 8690 8710
rect 7480 8680 7610 8690
rect 6300 8610 7310 8620
rect 6300 8470 6310 8610
rect 6860 8470 7310 8610
rect 6300 8460 7310 8470
rect 7770 8610 8790 8620
rect 7770 8470 8230 8610
rect 8780 8470 8790 8610
rect 7770 8460 8790 8470
rect 8830 8420 8980 8900
rect 9330 8850 10410 8860
rect 10540 9080 11620 9090
rect 11770 9040 11900 9050
rect 11760 8900 11770 9040
rect 11900 8900 11910 9040
rect 10540 8850 11620 8860
rect 9330 8710 9890 8850
rect 11060 8710 11620 8850
rect 9330 8700 10410 8710
rect 10540 8700 11620 8710
rect 10410 8680 10540 8690
rect 9230 8610 10240 8620
rect 9230 8470 9240 8610
rect 9790 8470 10240 8610
rect 9230 8460 10240 8470
rect 10700 8610 11720 8620
rect 10700 8470 11160 8610
rect 11710 8470 11720 8610
rect 10700 8460 11720 8470
rect 11760 8420 11910 8900
rect -20 8250 11910 8420
rect 1580 7300 3050 7460
rect 4420 7300 5890 7460
rect 7240 7300 8710 7460
rect 10150 7300 11620 7460
<< via2 >>
rect 1110 13380 2260 13820
rect 4040 13380 5190 13820
rect 6970 13380 8120 13820
rect 9900 13380 11050 13820
rect 380 11400 1010 12580
rect 2360 11400 2990 12580
rect 3310 11400 3940 12580
rect 5290 11400 5920 12580
rect 6240 11400 6870 12580
rect 8220 11400 8850 12580
rect 9170 11400 9800 12580
rect 11150 11400 11780 12580
rect 1110 10160 2260 10600
rect 4040 10160 5190 10600
rect 6970 10160 8120 10600
rect 9900 10160 11050 10600
rect 450 9330 1000 9470
rect 2370 9330 2920 9470
rect 1100 9090 1620 9230
rect 1620 9090 1750 9230
rect 1750 9090 2270 9230
rect 3380 9330 3930 9470
rect 5300 9330 5850 9470
rect 4030 9090 4550 9230
rect 4550 9090 4680 9230
rect 4680 9090 5200 9230
rect 1100 8710 1620 8850
rect 1620 8710 1750 8850
rect 1750 8710 2270 8850
rect 450 8470 1000 8610
rect 2370 8470 2920 8610
rect 6310 9330 6860 9470
rect 8230 9330 8780 9470
rect 6960 9090 7480 9230
rect 7480 9090 7610 9230
rect 7610 9090 8130 9230
rect 4030 8710 4550 8850
rect 4550 8710 4680 8850
rect 4680 8710 5200 8850
rect 3380 8470 3930 8610
rect 5300 8470 5850 8610
rect 9240 9330 9790 9470
rect 11160 9330 11710 9470
rect 9890 9090 10410 9230
rect 10410 9090 10540 9230
rect 10540 9090 11060 9230
rect 6960 8710 7480 8850
rect 7480 8710 7610 8850
rect 7610 8710 8130 8850
rect 6310 8470 6860 8610
rect 8230 8470 8780 8610
rect 9890 8710 10410 8850
rect 10410 8710 10540 8850
rect 10540 8710 11060 8850
rect 9240 8470 9790 8610
rect 11160 8470 11710 8610
<< metal3 >>
rect 210 13820 11950 14120
rect 210 13380 1110 13820
rect 2260 13380 4040 13820
rect 5190 13380 6970 13820
rect 8120 13380 9900 13820
rect 11050 13380 11950 13820
rect 210 12730 11950 13380
rect 370 12580 1020 12585
rect 370 11400 380 12580
rect 1010 11400 1020 12580
rect 370 11395 1020 11400
rect 440 9470 1010 11395
rect 1110 10605 2260 12730
rect 2350 12580 3000 12585
rect 2350 11400 2360 12580
rect 2350 11390 2380 11400
rect 2360 11360 2380 11390
rect 2990 11360 3000 12580
rect 3300 12580 3950 12585
rect 3300 11400 3310 12580
rect 3940 11400 3950 12580
rect 3300 11395 3950 11400
rect 1100 10600 2270 10605
rect 1100 10160 1110 10600
rect 2260 10160 2270 10600
rect 1100 10155 2270 10160
rect 440 9330 450 9470
rect 1000 9330 1010 9470
rect 440 8610 1010 9330
rect 2360 9470 2930 11360
rect 2360 9330 2370 9470
rect 2920 9330 2930 9470
rect 440 8470 450 8610
rect 1000 8470 1010 8610
rect 440 8460 1010 8470
rect 1090 9230 2280 9240
rect 1090 9090 1100 9230
rect 2270 9090 2280 9230
rect 1090 8850 2280 9090
rect 1090 8710 1100 8850
rect 2270 8710 2280 8850
rect 1090 8330 2280 8710
rect 2360 8610 2930 9330
rect 2360 8470 2370 8610
rect 2920 8470 2930 8610
rect 2360 8460 2930 8470
rect 3370 9470 3940 11395
rect 4040 10605 5190 12730
rect 5280 12580 5930 12585
rect 5280 11400 5290 12580
rect 5280 11395 5300 11400
rect 5290 11360 5300 11395
rect 5920 11360 5930 12580
rect 6230 12580 6880 12585
rect 6230 11400 6240 12580
rect 6870 11400 6880 12580
rect 6230 11395 6880 11400
rect 4030 10600 5200 10605
rect 4030 10160 4040 10600
rect 5190 10160 5200 10600
rect 4030 10155 5200 10160
rect 3370 9330 3380 9470
rect 3930 9330 3940 9470
rect 3370 8610 3940 9330
rect 5290 9470 5860 11360
rect 5290 9330 5300 9470
rect 5850 9330 5860 9470
rect 3370 8470 3380 8610
rect 3930 8470 3940 8610
rect 3370 8460 3940 8470
rect 4020 9230 5210 9240
rect 4020 9090 4030 9230
rect 5200 9090 5210 9230
rect 4020 8850 5210 9090
rect 4020 8710 4030 8850
rect 5200 8710 5210 8850
rect 4020 8330 5210 8710
rect 5290 8610 5860 9330
rect 5290 8470 5300 8610
rect 5850 8470 5860 8610
rect 5290 8460 5860 8470
rect 6300 9470 6870 11395
rect 6970 10605 8120 12730
rect 8210 12580 8860 12585
rect 8210 11360 8220 12580
rect 8850 11400 8860 12580
rect 8840 11395 8860 11400
rect 9160 12580 9810 12585
rect 9160 11400 9170 12580
rect 9800 11400 9810 12580
rect 9160 11395 9810 11400
rect 8840 11360 8850 11395
rect 6960 10600 8130 10605
rect 6960 10160 6970 10600
rect 8120 10160 8130 10600
rect 6960 10155 8130 10160
rect 6300 9330 6310 9470
rect 6860 9330 6870 9470
rect 6300 8610 6870 9330
rect 8220 9470 8790 11360
rect 8220 9330 8230 9470
rect 8780 9330 8790 9470
rect 6300 8470 6310 8610
rect 6860 8470 6870 8610
rect 6300 8460 6870 8470
rect 6950 9230 8140 9240
rect 6950 9090 6960 9230
rect 8130 9090 8140 9230
rect 6950 8850 8140 9090
rect 6950 8710 6960 8850
rect 8130 8710 8140 8850
rect 6950 8330 8140 8710
rect 8220 8610 8790 9330
rect 8220 8470 8230 8610
rect 8780 8470 8790 8610
rect 8220 8460 8790 8470
rect 9230 9470 9800 11395
rect 9900 10605 11050 12730
rect 11140 12580 11790 12585
rect 11140 11400 11150 12580
rect 11140 11395 11160 11400
rect 11150 11360 11160 11395
rect 11780 11360 11790 12580
rect 9890 10600 11060 10605
rect 9890 10160 9900 10600
rect 11050 10160 11060 10600
rect 9890 10155 11060 10160
rect 9230 9330 9240 9470
rect 9790 9330 9800 9470
rect 9230 8610 9800 9330
rect 11150 9470 11720 11360
rect 11150 9330 11160 9470
rect 11710 9330 11720 9470
rect 9230 8470 9240 8610
rect 9790 8470 9800 8610
rect 9230 8460 9800 8470
rect 9880 9230 11070 9240
rect 9880 9090 9890 9230
rect 11060 9090 11070 9230
rect 9880 8850 11070 9090
rect 9880 8710 9890 8850
rect 11060 8710 11070 8850
rect 9880 8330 11070 8710
rect 11150 8610 11720 9330
rect 11150 8470 11160 8610
rect 11710 8470 11720 8610
rect 11150 8460 11720 8470
rect 960 8130 13100 8330
rect 950 7840 13100 8130
rect 950 7560 13090 7840
rect 970 140 1880 450
rect 3820 140 4730 460
rect 6670 140 7580 450
rect 9520 140 10430 450
rect 12370 140 13280 450
rect -20 -880 14220 140
<< via3 >>
rect 380 12040 1000 12560
rect 2380 11400 2990 11880
rect 2380 11360 2990 11400
rect 3320 12040 3940 12560
rect 5300 11400 5920 11880
rect 5300 11360 5920 11400
rect 6240 12040 6860 12560
rect 8220 11400 8840 11880
rect 8220 11360 8840 11400
rect 9180 12040 9800 12560
rect 11160 11400 11780 11880
rect 11160 11360 11780 11400
<< metal4 >>
rect 360 12560 11960 12580
rect 360 12040 380 12560
rect 1000 12040 3320 12560
rect 3940 12040 6240 12560
rect 6860 12040 9180 12560
rect 9800 12040 11960 12560
rect 360 12020 11960 12040
rect 360 11880 11960 11900
rect 360 11360 2380 11880
rect 2990 11360 5300 11880
rect 5920 11360 8220 11880
rect 8840 11360 11160 11880
rect 11780 11360 11960 11880
rect 360 11340 11960 11360
use outd_cmirror_64t#1  outd_cmirror_64t_0
timestamp 1646921651
transform 1 0 -30 0 1 76
box 0 -76 2862 7840
use outd_cmirror_64t#1  outd_cmirror_64t_1
timestamp 1646921651
transform 1 0 2820 0 1 76
box 0 -76 2862 7840
use outd_cmirror_64t#1  outd_cmirror_64t_2
timestamp 1646921651
transform 1 0 5670 0 1 76
box 0 -76 2862 7840
use outd_cmirror_64t#1  outd_cmirror_64t_3
timestamp 1646921651
transform 1 0 8520 0 1 76
box 0 -76 2862 7840
use outd_cmirror_64t#1  outd_cmirror_64t_4
timestamp 1646921651
transform 1 0 11370 0 1 76
box 0 -76 2862 7840
use outd_diffamp#1  outd_diffamp_0
timestamp 1646921651
transform 1 0 300 0 1 320
box 0 7930 2768 9368
use outd_diffamp#1  outd_diffamp_1
timestamp 1646921651
transform 1 0 3230 0 1 320
box 0 7930 2768 9368
use outd_diffamp#1  outd_diffamp_2
timestamp 1646921651
transform 1 0 6160 0 1 320
box 0 7930 2768 9368
use outd_diffamp#1  outd_diffamp_3
timestamp 1646921651
transform 1 0 9090 0 1 320
box 0 7930 2768 9368
use sky130_fd_pr__res_high_po_5p73_PA2QZX  sky130_fd_pr__res_high_po_5p73_PA2QZX_0
timestamp 1646921651
transform 1 0 951 0 1 10998
box -739 -998 739 998
use sky130_fd_pr__res_high_po_5p73_PA2QZX  sky130_fd_pr__res_high_po_5p73_PA2QZX_1
timestamp 1646921651
transform 1 0 2419 0 1 10998
box -739 -998 739 998
use sky130_fd_pr__res_high_po_5p73_PA2QZX  sky130_fd_pr__res_high_po_5p73_PA2QZX_2
timestamp 1646921651
transform 1 0 951 0 1 12978
box -739 -998 739 998
use sky130_fd_pr__res_high_po_5p73_PA2QZX  sky130_fd_pr__res_high_po_5p73_PA2QZX_3
timestamp 1646921651
transform 1 0 2419 0 1 12978
box -739 -998 739 998
use sky130_fd_pr__res_high_po_5p73_PA2QZX  sky130_fd_pr__res_high_po_5p73_PA2QZX_4
timestamp 1646921651
transform 1 0 5349 0 1 10998
box -739 -998 739 998
use sky130_fd_pr__res_high_po_5p73_PA2QZX  sky130_fd_pr__res_high_po_5p73_PA2QZX_5
timestamp 1646921651
transform 1 0 3881 0 1 10998
box -739 -998 739 998
use sky130_fd_pr__res_high_po_5p73_PA2QZX  sky130_fd_pr__res_high_po_5p73_PA2QZX_6
timestamp 1646921651
transform 1 0 3881 0 1 12978
box -739 -998 739 998
use sky130_fd_pr__res_high_po_5p73_PA2QZX  sky130_fd_pr__res_high_po_5p73_PA2QZX_7
timestamp 1646921651
transform 1 0 5349 0 1 12978
box -739 -998 739 998
use sky130_fd_pr__res_high_po_5p73_PA2QZX  sky130_fd_pr__res_high_po_5p73_PA2QZX_8
timestamp 1646921651
transform 1 0 8279 0 1 10998
box -739 -998 739 998
use sky130_fd_pr__res_high_po_5p73_PA2QZX  sky130_fd_pr__res_high_po_5p73_PA2QZX_9
timestamp 1646921651
transform 1 0 6811 0 1 10998
box -739 -998 739 998
use sky130_fd_pr__res_high_po_5p73_PA2QZX  sky130_fd_pr__res_high_po_5p73_PA2QZX_10
timestamp 1646921651
transform 1 0 6811 0 1 12978
box -739 -998 739 998
use sky130_fd_pr__res_high_po_5p73_PA2QZX  sky130_fd_pr__res_high_po_5p73_PA2QZX_11
timestamp 1646921651
transform 1 0 8279 0 1 12978
box -739 -998 739 998
use sky130_fd_pr__res_high_po_5p73_PA2QZX  sky130_fd_pr__res_high_po_5p73_PA2QZX_12
timestamp 1646921651
transform 1 0 11209 0 1 10998
box -739 -998 739 998
use sky130_fd_pr__res_high_po_5p73_PA2QZX  sky130_fd_pr__res_high_po_5p73_PA2QZX_13
timestamp 1646921651
transform 1 0 9741 0 1 10998
box -739 -998 739 998
use sky130_fd_pr__res_high_po_5p73_PA2QZX  sky130_fd_pr__res_high_po_5p73_PA2QZX_14
timestamp 1646921651
transform 1 0 9741 0 1 12978
box -739 -998 739 998
use sky130_fd_pr__res_high_po_5p73_PA2QZX  sky130_fd_pr__res_high_po_5p73_PA2QZX_15
timestamp 1646921651
transform 1 0 11209 0 1 12978
box -739 -998 739 998
<< labels >>
rlabel metal3 2384 7668 2640 7832 1 cmirror_out
rlabel metal3 240 -442 496 -278 1 VN
<< end >>
