magic
tech sky130A
magscale 1 2
timestamp 1647254192
<< pwell >>
rect -941 -410 941 410
<< nmos >>
rect -745 -200 -545 200
rect -487 -200 -287 200
rect -229 -200 -29 200
rect 29 -200 229 200
rect 287 -200 487 200
rect 545 -200 745 200
<< ndiff >>
rect -803 188 -745 200
rect -803 -188 -791 188
rect -757 -188 -745 188
rect -803 -200 -745 -188
rect -545 188 -487 200
rect -545 -188 -533 188
rect -499 -188 -487 188
rect -545 -200 -487 -188
rect -287 188 -229 200
rect -287 -188 -275 188
rect -241 -188 -229 188
rect -287 -200 -229 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 229 188 287 200
rect 229 -188 241 188
rect 275 -188 287 188
rect 229 -200 287 -188
rect 487 188 545 200
rect 487 -188 499 188
rect 533 -188 545 188
rect 487 -200 545 -188
rect 745 188 803 200
rect 745 -188 757 188
rect 791 -188 803 188
rect 745 -200 803 -188
<< ndiffc >>
rect -791 -188 -757 188
rect -533 -188 -499 188
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
rect 499 -188 533 188
rect 757 -188 791 188
<< psubdiff >>
rect -905 340 -809 374
rect 809 340 905 374
rect -905 278 -871 340
rect 871 278 905 340
rect -905 -340 -871 -278
rect 871 -340 905 -278
rect -905 -374 -809 -340
rect 809 -374 905 -340
<< psubdiffcont >>
rect -809 340 809 374
rect -905 -278 -871 278
rect 871 -278 905 278
rect -809 -374 809 -340
<< poly >>
rect -745 272 -545 288
rect -745 238 -729 272
rect -561 238 -545 272
rect -745 200 -545 238
rect -487 272 -287 288
rect -487 238 -471 272
rect -303 238 -287 272
rect -487 200 -287 238
rect -229 272 -29 288
rect -229 238 -213 272
rect -45 238 -29 272
rect -229 200 -29 238
rect 29 272 229 288
rect 29 238 45 272
rect 213 238 229 272
rect 29 200 229 238
rect 287 272 487 288
rect 287 238 303 272
rect 471 238 487 272
rect 287 200 487 238
rect 545 272 745 288
rect 545 238 561 272
rect 729 238 745 272
rect 545 200 745 238
rect -745 -238 -545 -200
rect -745 -272 -729 -238
rect -561 -272 -545 -238
rect -745 -288 -545 -272
rect -487 -238 -287 -200
rect -487 -272 -471 -238
rect -303 -272 -287 -238
rect -487 -288 -287 -272
rect -229 -238 -29 -200
rect -229 -272 -213 -238
rect -45 -272 -29 -238
rect -229 -288 -29 -272
rect 29 -238 229 -200
rect 29 -272 45 -238
rect 213 -272 229 -238
rect 29 -288 229 -272
rect 287 -238 487 -200
rect 287 -272 303 -238
rect 471 -272 487 -238
rect 287 -288 487 -272
rect 545 -238 745 -200
rect 545 -272 561 -238
rect 729 -272 745 -238
rect 545 -288 745 -272
<< polycont >>
rect -729 238 -561 272
rect -471 238 -303 272
rect -213 238 -45 272
rect 45 238 213 272
rect 303 238 471 272
rect 561 238 729 272
rect -729 -272 -561 -238
rect -471 -272 -303 -238
rect -213 -272 -45 -238
rect 45 -272 213 -238
rect 303 -272 471 -238
rect 561 -272 729 -238
<< locali >>
rect -905 340 -809 374
rect 809 340 905 374
rect -905 278 -871 340
rect 871 278 905 340
rect -745 238 -729 272
rect -561 238 -545 272
rect -487 238 -471 272
rect -303 238 -287 272
rect -229 238 -213 272
rect -45 238 -29 272
rect 29 238 45 272
rect 213 238 229 272
rect 287 238 303 272
rect 471 238 487 272
rect 545 238 561 272
rect 729 238 745 272
rect -791 188 -757 204
rect -791 -204 -757 -188
rect -533 188 -499 204
rect -533 -204 -499 -188
rect -275 188 -241 204
rect -275 -204 -241 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 241 188 275 204
rect 241 -204 275 -188
rect 499 188 533 204
rect 499 -204 533 -188
rect 757 188 791 204
rect 757 -204 791 -188
rect -745 -272 -729 -238
rect -561 -272 -545 -238
rect -487 -272 -471 -238
rect -303 -272 -287 -238
rect -229 -272 -213 -238
rect -45 -272 -29 -238
rect 29 -272 45 -238
rect 213 -272 229 -238
rect 287 -272 303 -238
rect 471 -272 487 -238
rect 545 -272 561 -238
rect 729 -272 745 -238
rect -905 -340 -871 -278
rect 871 -340 905 -278
rect -905 -374 -809 -340
rect 809 -374 905 -340
<< viali >>
rect -729 238 -561 272
rect -471 238 -303 272
rect -213 238 -45 272
rect 45 238 213 272
rect 303 238 471 272
rect 561 238 729 272
rect -791 -188 -757 188
rect -533 -188 -499 188
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
rect 499 -188 533 188
rect 757 -188 791 188
rect -729 -272 -561 -238
rect -471 -272 -303 -238
rect -213 -272 -45 -238
rect 45 -272 213 -238
rect 303 -272 471 -238
rect 561 -272 729 -238
<< metal1 >>
rect -741 272 -549 278
rect -741 238 -729 272
rect -561 238 -549 272
rect -741 232 -549 238
rect -483 272 -291 278
rect -483 238 -471 272
rect -303 238 -291 272
rect -483 232 -291 238
rect -225 272 -33 278
rect -225 238 -213 272
rect -45 238 -33 272
rect -225 232 -33 238
rect 33 272 225 278
rect 33 238 45 272
rect 213 238 225 272
rect 33 232 225 238
rect 291 272 483 278
rect 291 238 303 272
rect 471 238 483 272
rect 291 232 483 238
rect 549 272 741 278
rect 549 238 561 272
rect 729 238 741 272
rect 549 232 741 238
rect -797 188 -751 200
rect -797 -188 -791 188
rect -757 -188 -751 188
rect -797 -200 -751 -188
rect -539 188 -493 200
rect -539 -188 -533 188
rect -499 -188 -493 188
rect -539 -200 -493 -188
rect -281 188 -235 200
rect -281 -188 -275 188
rect -241 -188 -235 188
rect -281 -200 -235 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 235 188 281 200
rect 235 -188 241 188
rect 275 -188 281 188
rect 235 -200 281 -188
rect 493 188 539 200
rect 493 -188 499 188
rect 533 -188 539 188
rect 493 -200 539 -188
rect 751 188 797 200
rect 751 -188 757 188
rect 791 -188 797 188
rect 751 -200 797 -188
rect -741 -238 -549 -232
rect -741 -272 -729 -238
rect -561 -272 -549 -238
rect -741 -278 -549 -272
rect -483 -238 -291 -232
rect -483 -272 -471 -238
rect -303 -272 -291 -238
rect -483 -278 -291 -272
rect -225 -238 -33 -232
rect -225 -272 -213 -238
rect -45 -272 -33 -238
rect -225 -278 -33 -272
rect 33 -238 225 -232
rect 33 -272 45 -238
rect 213 -272 225 -238
rect 33 -278 225 -272
rect 291 -238 483 -232
rect 291 -272 303 -238
rect 471 -272 483 -238
rect 291 -278 483 -272
rect 549 -238 741 -232
rect 549 -272 561 -238
rect 729 -272 741 -238
rect 549 -278 741 -272
<< properties >>
string FIXED_BBOX -888 -357 888 357
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 1 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
