* SPICE3 file created from tia_one_tia.ext - technology: sky130A

X0 tia_cur_mirror_0/m1_71_130# tia_cur_mirror_0/a_122_42# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1 tia_cur_mirror_0/m1_71_130# tia_cur_mirror_0/a_122_42# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2 m1_1540_1550# tia_cur_mirror_0/a_122_42# tia_cur_mirror_0/m1_71_130# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3 m1_1540_1550# tia_cur_mirror_0/a_122_42# tia_cur_mirror_0/m1_71_130# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4 tia_cur_mirror_0/m1_71_130# tia_cur_mirror_0/a_122_42# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5 tia_cur_mirror_0/m1_71_130# tia_cur_mirror_0/a_122_42# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6 tia_cur_mirror_0/m1_71_130# tia_cur_mirror_0/a_122_42# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7 m1_1540_1550# tia_cur_mirror_0/a_122_42# tia_cur_mirror_0/m1_71_130# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8 m1_1540_1550# tia_cur_mirror_0/a_122_42# tia_cur_mirror_0/m1_71_130# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9 m1_1540_1550# tia_cur_mirror_0/a_122_42# tia_cur_mirror_0/m1_71_130# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10 m1_1540_1550# tia_cur_mirror_0/a_122_42# tia_cur_mirror_0/m1_71_130# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11 tia_cur_mirror_0/m1_71_130# tia_cur_mirror_0/a_122_42# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12 VSUBS tia_cur_mirror_0/a_122_42# tia_cur_mirror_0/m1_71_130# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13 tia_cur_mirror_0/m1_71_130# tia_cur_mirror_0/a_122_42# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14 tia_cur_mirror_0/m1_71_130# tia_cur_mirror_0/a_122_42# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15 VSUBS tia_cur_mirror_0/a_122_42# tia_cur_mirror_0/m1_71_130# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X16 tia_cur_mirror_0/m1_71_130# tia_cur_mirror_0/a_122_42# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X17 VSUBS tia_cur_mirror_0/a_122_42# tia_cur_mirror_0/m1_71_130# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X18 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X19 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X20 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X21 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X22 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X23 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X24 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X25 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X26 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X27 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X28 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X29 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X30 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X31 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X32 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X33 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X34 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X35 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X36 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X37 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X38 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X39 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X40 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X41 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X42 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X43 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X44 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X45 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X46 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X47 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X48 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X49 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X50 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X51 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X52 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X53 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X54 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X55 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X56 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X57 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X58 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X59 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X60 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X61 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X62 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X63 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X64 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X65 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X66 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X67 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X68 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X69 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X70 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X71 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X72 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X73 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X74 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X75 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X76 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X77 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X78 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X79 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X80 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X81 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X82 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X83 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X84 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X85 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X86 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X87 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X88 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X89 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X90 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X91 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X92 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X93 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X94 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X95 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X96 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X97 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X98 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X99 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X100 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X101 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X102 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X103 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X104 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X105 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X106 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X107 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X108 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X109 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X110 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X111 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X112 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X113 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X114 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X115 m1_1540_1550# w_1686_386# m2_n1710_n500# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X116 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X117 m2_n1710_n500# w_1686_386# m1_1540_1550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X118 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X119 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X120 m1_1540_1550# w_1686_386# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X121 m1_1540_1550# w_1686_386# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X122 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X123 m1_1540_1550# w_1686_386# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X124 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X125 m1_1540_1550# w_1686_386# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X126 m1_1540_1550# w_1686_386# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X127 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X128 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X129 m1_1540_1550# w_1686_386# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X130 m1_1540_1550# w_1686_386# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X131 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X132 m1_1540_1550# w_1686_386# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X133 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X134 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X135 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X136 m1_1540_1550# w_1686_386# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X137 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X138 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X139 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X140 m1_1540_1550# w_1686_386# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X141 m1_1540_1550# w_1686_386# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X142 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X143 m1_1540_1550# w_1686_386# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X144 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X145 m1_1540_1550# w_1686_386# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X146 m1_1540_1550# w_1686_386# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X147 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X148 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X149 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X150 m1_1540_1550# w_1686_386# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X151 m1_1540_1550# w_1686_386# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X152 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X153 m1_1540_1550# w_1686_386# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X154 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X155 m1_1540_1550# w_1686_386# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X156 m1_1540_1550# w_1686_386# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X157 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X158 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X159 m1_1540_1550# w_1686_386# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X160 m1_1540_1550# w_1686_386# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X161 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X162 m1_1540_1550# w_1686_386# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X163 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X164 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X165 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X166 m1_1540_1550# w_1686_386# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X167 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X168 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X169 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X170 m1_1540_1550# w_1686_386# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X171 m1_1540_1550# w_1686_386# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X172 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X173 m1_1540_1550# w_1686_386# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X174 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X175 m1_1540_1550# w_1686_386# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X176 m1_1540_1550# w_1686_386# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X177 w_1650_2620# w_1686_386# m1_1540_1550# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X178 w_1650_2620# sky130_fd_pr__cap_mim_m3_2_ZWVPUJ_0/m4_n2851_n1900# sky130_fd_pr__cap_mim_m3_2 l=1.8e+07u w=2.5e+07u
X179 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X180 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X181 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X182 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X183 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X184 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X185 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X186 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X187 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X188 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X189 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X190 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X191 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X192 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X193 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X194 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X195 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X196 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X197 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X198 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X199 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X200 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X201 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X202 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X203 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X204 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X205 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X206 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X207 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X208 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X209 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X210 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X211 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X212 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X213 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X214 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X215 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X216 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X217 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X218 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X219 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X220 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X221 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X222 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X223 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X224 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X225 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X226 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X227 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X228 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X229 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X230 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X231 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X232 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X233 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X234 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X235 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X236 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X237 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X238 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X239 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X240 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X241 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X242 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X243 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X244 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X245 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X246 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X247 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X248 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X249 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X250 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X251 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X252 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X253 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X254 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X255 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X256 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X257 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X258 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X259 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X260 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X261 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X262 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X263 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X264 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X265 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X266 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X267 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X268 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X269 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X270 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X271 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X272 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X273 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X274 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X275 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X276 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X277 VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X278 m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X279 m2_1800_2380# m1_1850_2290# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X280 m2_1800_2380# m1_1850_2290# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X281 w_1650_2620# m1_1850_2290# m2_1800_2380# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X282 w_1650_2620# m1_1850_2290# m2_1800_2380# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X283 m2_1800_2380# m1_1850_2290# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X284 m2_1800_2380# m1_1850_2290# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X285 m2_1800_2380# m1_1850_2290# w_1650_2620# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X286 w_1650_2620# m1_1850_2290# m2_1800_2380# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X287 w_1650_2620# m1_1850_2290# m2_1800_2380# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X288 w_1650_2620# m1_1850_2290# m2_1800_2380# w_1650_2620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X289 w_1686_386# m1_1540_1550# m2_1800_2380# w_1686_386# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X290 w_1686_386# m1_1540_1550# m2_1800_2380# w_1686_386# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X291 m2_1800_2380# m1_1540_1550# w_1686_386# w_1686_386# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X292 m2_1800_2380# m1_1540_1550# w_1686_386# w_1686_386# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X293 w_1686_386# m1_1540_1550# m2_1800_2380# w_1686_386# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X294 m2_1800_2380# m1_1540_1550# w_1686_386# w_1686_386# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X295 w_1686_386# m1_1540_1550# m2_1800_2380# w_1686_386# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X296 w_1686_386# m1_1540_1550# m2_1800_2380# w_1686_386# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X297 w_1686_386# m1_1540_1550# m2_1800_2380# w_1686_386# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X298 m2_1800_2380# m1_1540_1550# w_1686_386# w_1686_386# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X299 w_1686_386# m1_1540_1550# m2_1800_2380# w_1686_386# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X300 w_1686_386# m1_1540_1550# m2_1800_2380# w_1686_386# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X301 w_1686_386# m1_1540_1550# m2_1800_2380# w_1686_386# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X302 m2_1800_2380# m1_1540_1550# w_1686_386# w_1686_386# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X303 m2_1800_2380# m1_1540_1550# w_1686_386# w_1686_386# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X304 m2_1800_2380# m1_1540_1550# w_1686_386# w_1686_386# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X305 w_1686_386# m1_1540_1550# m2_1800_2380# w_1686_386# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X306 w_1686_386# m1_1540_1550# m2_1800_2380# w_1686_386# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X307 m2_1800_2380# m1_1540_1550# w_1686_386# w_1686_386# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X308 m2_1800_2380# m1_1540_1550# w_1686_386# w_1686_386# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X309 w_1686_386# m1_1540_1550# m2_1800_2380# w_1686_386# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X310 w_1686_386# m1_1540_1550# m2_1800_2380# w_1686_386# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X311 w_1686_386# m1_1540_1550# m2_1800_2380# w_1686_386# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X312 m2_1800_2380# m1_1540_1550# w_1686_386# w_1686_386# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X313 m2_1800_2380# m1_1540_1550# w_1686_386# w_1686_386# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X314 w_1686_386# m1_1540_1550# m2_1800_2380# w_1686_386# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X315 m2_1800_2380# m1_1540_1550# w_1686_386# w_1686_386# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X316 w_1686_386# m1_1540_1550# m2_1800_2380# w_1686_386# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X317 m2_1800_2380# m1_1540_1550# w_1686_386# w_1686_386# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X318 m2_1800_2380# m1_1540_1550# w_1686_386# w_1686_386# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
