magic
tech sky130A
timestamp 1647254192
<< nwell >>
rect -1005 640 -980 985
<< pwell >>
rect -4320 160 -4220 510
rect -3910 155 -3810 505
rect -3505 150 -3405 500
rect -3095 150 -2995 500
rect -2690 150 -2590 500
rect -2280 150 -2180 500
rect -1870 150 -1770 500
rect -1460 150 -1360 500
rect -1055 150 -955 500
rect -645 150 -555 550
<< locali >>
rect -4715 1055 -555 1095
rect -4715 550 -4680 1055
rect -4565 935 -4290 940
rect -4565 670 -4560 935
rect -4295 670 -4290 935
rect -4565 665 -4290 670
rect -4170 935 -3890 940
rect -4170 670 -4160 935
rect -3895 670 -3890 935
rect -4170 665 -3890 670
rect -3770 935 -3490 940
rect -3770 670 -3765 935
rect -3495 670 -3490 935
rect -3770 665 -3490 670
rect -3370 935 -3095 940
rect -3370 670 -3365 935
rect -3100 670 -3095 935
rect -3370 665 -3095 670
rect -2975 935 -2695 940
rect -2975 670 -2970 935
rect -2700 670 -2695 935
rect -2975 665 -2695 670
rect -2575 935 -2300 940
rect -2575 670 -2570 935
rect -2305 670 -2300 935
rect -2575 665 -2300 670
rect -2180 935 -1900 940
rect -2180 670 -2175 935
rect -1905 670 -1900 935
rect -2180 665 -1900 670
rect -1780 935 -1500 940
rect -1780 670 -1775 935
rect -1505 670 -1500 935
rect -1780 665 -1500 670
rect -1385 670 -1375 940
rect -1105 670 -1100 940
rect -1385 665 -1100 670
rect -985 670 -980 940
rect -710 670 -705 940
rect -985 665 -705 670
rect -590 550 -555 1055
rect -560 150 -555 550
<< viali >>
rect -4600 940 -665 985
rect -4600 665 -4565 940
rect -4290 665 -4170 940
rect -3890 665 -3770 940
rect -3490 665 -3370 940
rect -3095 665 -2975 940
rect -2695 665 -2575 940
rect -2300 665 -2180 940
rect -1900 665 -1780 940
rect -1500 665 -1385 940
rect -1100 665 -985 940
rect -705 665 -665 940
rect -4600 625 -665 665
rect -4715 485 -560 550
rect -4715 190 -4620 485
rect -4325 190 -4215 485
rect -3915 190 -3805 485
rect -3510 190 -3400 485
rect -3100 190 -2990 485
rect -2695 190 -2585 485
rect -2285 190 -2175 485
rect -1875 190 -1765 485
rect -1470 190 -1360 485
rect -1060 190 -950 485
rect -655 190 -560 485
rect -4715 150 -560 190
<< metal1 >>
rect -4605 988 -660 1095
rect -4606 985 -659 988
rect -4606 937 -4600 985
rect -4603 668 -4600 937
rect -4606 625 -4600 668
rect -4565 937 -4290 940
rect -4565 668 -4562 937
rect -4530 710 -4525 895
rect -4335 710 -4330 895
rect -4293 668 -4290 937
rect -4565 665 -4290 668
rect -4170 937 -3890 940
rect -4170 668 -4167 937
rect -4130 710 -4125 895
rect -3935 710 -3930 895
rect -3893 668 -3890 937
rect -4170 665 -3890 668
rect -3770 937 -3490 940
rect -3770 668 -3767 937
rect -3730 710 -3725 895
rect -3535 710 -3530 895
rect -3493 668 -3490 937
rect -3770 665 -3490 668
rect -3370 937 -3095 940
rect -3370 668 -3367 937
rect -3335 710 -3330 895
rect -3140 710 -3135 895
rect -3098 668 -3095 937
rect -3370 665 -3095 668
rect -2975 937 -2695 940
rect -2975 668 -2972 937
rect -2935 710 -2930 895
rect -2740 710 -2735 895
rect -2698 668 -2695 937
rect -2975 665 -2695 668
rect -2575 937 -2300 940
rect -2575 668 -2572 937
rect -2540 710 -2535 895
rect -2345 710 -2340 895
rect -2303 668 -2300 937
rect -2575 665 -2300 668
rect -2180 937 -1900 940
rect -2180 668 -2177 937
rect -2140 710 -2135 895
rect -1945 710 -1940 895
rect -1903 668 -1900 937
rect -2180 665 -1900 668
rect -1780 937 -1500 940
rect -1780 668 -1777 937
rect -1740 710 -1735 895
rect -1545 710 -1540 895
rect -1503 668 -1500 937
rect -1780 665 -1500 668
rect -1385 937 -1100 940
rect -1385 668 -1382 937
rect -1340 710 -1335 895
rect -1150 710 -1145 895
rect -1103 668 -1100 937
rect -1385 665 -1100 668
rect -985 937 -705 940
rect -985 668 -982 937
rect -940 710 -935 895
rect -750 710 -745 895
rect -708 668 -705 937
rect -985 665 -705 668
rect -665 937 -659 985
rect -665 668 -662 937
rect -665 625 -659 668
rect -4606 622 -659 625
rect -4603 619 -4562 622
rect -4293 619 -4167 622
rect -3893 619 -3767 622
rect -3493 619 -3367 622
rect -3098 619 -2972 622
rect -2698 619 -2572 622
rect -2303 619 -2177 622
rect -1903 619 -1777 622
rect -1503 619 -1382 622
rect -1103 619 -982 622
rect -708 619 -662 622
rect -4718 553 -4617 556
rect -4328 553 -4212 556
rect -3918 553 -3802 556
rect -3513 553 -3397 556
rect -3103 553 -2987 556
rect -2698 553 -2582 556
rect -2288 553 -2172 556
rect -1878 553 -1762 556
rect -1473 553 -1357 556
rect -1063 553 -947 556
rect -658 553 -557 556
rect -4721 550 -554 553
rect -4721 482 -4715 550
rect -4718 193 -4715 482
rect -4721 150 -4715 193
rect -4620 482 -4325 485
rect -4620 193 -4617 482
rect -4570 245 -4565 425
rect -4385 245 -4380 425
rect -4328 193 -4325 482
rect -4620 190 -4325 193
rect -4215 482 -3915 485
rect -4215 193 -4212 482
rect -4160 245 -4155 425
rect -3975 245 -3970 425
rect -3918 193 -3915 482
rect -4215 190 -3915 193
rect -3805 482 -3510 485
rect -3805 193 -3802 482
rect -3755 245 -3750 430
rect -3565 245 -3560 430
rect -3513 193 -3510 482
rect -3805 190 -3510 193
rect -3400 482 -3100 485
rect -3400 193 -3397 482
rect -3345 245 -3340 430
rect -3155 245 -3150 430
rect -3103 193 -3100 482
rect -3400 190 -3100 193
rect -2990 482 -2695 485
rect -2990 193 -2987 482
rect -2940 245 -2935 430
rect -2750 245 -2745 430
rect -2698 193 -2695 482
rect -2990 190 -2695 193
rect -2585 482 -2285 485
rect -2585 193 -2582 482
rect -2530 245 -2525 430
rect -2340 245 -2335 430
rect -2288 193 -2285 482
rect -2585 190 -2285 193
rect -2175 482 -1875 485
rect -2175 193 -2172 482
rect -2125 245 -2120 430
rect -1935 245 -1930 430
rect -1878 193 -1875 482
rect -2175 190 -1875 193
rect -1765 482 -1470 485
rect -1765 193 -1762 482
rect -1715 245 -1710 430
rect -1525 245 -1520 430
rect -1473 193 -1470 482
rect -1765 190 -1470 193
rect -1360 482 -1060 485
rect -1360 193 -1357 482
rect -1305 245 -1300 430
rect -1115 245 -1110 430
rect -1063 193 -1060 482
rect -1360 190 -1060 193
rect -950 482 -655 485
rect -950 193 -947 482
rect -900 245 -895 430
rect -710 245 -705 430
rect -658 193 -655 482
rect -950 190 -655 193
rect -560 482 -554 550
rect -560 193 -557 482
rect -560 150 -554 193
rect -4721 147 -554 150
rect -4718 144 -4617 147
rect -4328 144 -4212 147
rect -3918 144 -3802 147
rect -3513 144 -3397 147
rect -3103 144 -2987 147
rect -2698 144 -2582 147
rect -2288 144 -2172 147
rect -1878 144 -1762 147
rect -1473 144 -1357 147
rect -1063 144 -947 147
rect -658 144 -557 147
<< via1 >>
rect -4525 710 -4335 895
rect -4125 710 -3935 895
rect -3725 710 -3535 895
rect -3330 710 -3140 895
rect -2930 710 -2740 895
rect -2535 710 -2345 895
rect -2135 710 -1945 895
rect -1735 710 -1545 895
rect -1335 710 -1150 895
rect -935 710 -750 895
rect -4565 245 -4385 425
rect -4155 245 -3975 425
rect -3750 245 -3565 430
rect -3340 245 -3155 430
rect -2935 245 -2750 430
rect -2525 245 -2340 430
rect -2120 245 -1935 430
rect -1710 245 -1525 430
rect -1300 245 -1115 430
rect -895 245 -710 430
<< metal2 >>
rect -4570 895 -705 905
rect -4570 710 -4525 895
rect -4335 710 -4125 895
rect -3935 710 -3725 895
rect -3535 710 -3330 895
rect -3140 710 -2930 895
rect -2740 710 -2535 895
rect -2345 710 -2135 895
rect -1945 710 -1735 895
rect -1545 710 -1335 895
rect -1150 710 -935 895
rect -750 710 -705 895
rect -4570 430 -705 710
rect -4570 425 -3750 430
rect -4570 245 -4565 425
rect -4385 245 -4155 425
rect -3975 245 -3750 425
rect -3565 245 -3340 430
rect -3155 245 -2935 430
rect -2750 245 -2525 430
rect -2340 245 -2120 430
rect -1935 245 -1710 430
rect -1525 245 -1300 430
rect -1115 245 -895 430
rect -710 245 -705 430
rect -4570 240 -705 245
use sky130_fd_pr__diode_pd2nw_11v0_33C8ED  sky130_fd_pr__diode_pd2nw_11v0_33C8ED_0
timestamp 1647254192
transform 1 0 -2635 0 1 804
box -2080 -289 2080 289
use sky130_fd_pr__diode_pw2nd_11v0_T9UBGD  sky130_fd_pr__diode_pw2nd_11v0_T9UBGD_0
timestamp 1647254192
transform 1 0 -2638 0 1 336
box -2022 -186 2022 186
<< end >>
