magic
tech sky130A
magscale 1 2
timestamp 1647254192
<< locali >>
rect 0 2200 2040 2280
rect 0 60 60 2200
rect 380 1840 480 2200
rect 1980 2020 2040 2200
rect 1880 1840 2040 2020
rect 360 320 480 1840
rect 1980 420 2040 1840
rect 380 60 480 320
rect 1880 240 2040 420
rect 1980 60 2040 240
rect 0 0 2040 60
<< metal1 >>
rect 100 2120 1860 2180
rect 100 2100 1850 2120
rect 180 2090 260 2100
rect 110 1260 120 1460
rect 180 1260 190 1460
rect 250 1260 260 1460
rect 320 1260 330 1460
rect 360 1220 480 2100
rect 810 1840 820 2040
rect 880 1840 890 2040
rect 1330 1840 1340 2040
rect 1400 1840 1410 2040
rect 1830 1840 1840 2040
rect 1920 1840 1930 2040
rect 550 1260 560 1460
rect 620 1260 630 1460
rect 1070 1260 1080 1460
rect 1140 1260 1150 1460
rect 1590 1260 1600 1460
rect 1660 1260 1670 1460
rect 0 1060 1880 1220
rect 110 820 120 1020
rect 180 820 190 1020
rect 250 820 260 1020
rect 320 820 330 1020
rect 360 180 480 1060
rect 550 820 560 1020
rect 620 820 630 1020
rect 1070 820 1080 1020
rect 1140 820 1150 1020
rect 1590 820 1600 1020
rect 1660 820 1670 1020
rect 810 220 820 420
rect 880 220 890 420
rect 1330 220 1340 420
rect 1400 220 1410 420
rect 1830 220 1840 420
rect 1920 220 1930 420
rect 100 160 1850 180
rect 100 100 1860 160
<< via1 >>
rect 120 1260 180 1460
rect 260 1260 320 1460
rect 820 1840 880 2040
rect 1340 1840 1400 2040
rect 1840 1840 1920 2040
rect 560 1260 620 1460
rect 1080 1260 1140 1460
rect 1600 1260 1660 1460
rect 120 820 180 1020
rect 260 820 320 1020
rect 560 820 620 1020
rect 1080 820 1140 1020
rect 1600 820 1660 1020
rect 820 220 880 420
rect 1340 220 1400 420
rect 1840 220 1920 420
<< metal2 >>
rect 820 2040 880 2050
rect 1340 2040 1400 2050
rect 1840 2040 1920 2050
rect 880 1840 1340 2040
rect 1400 1840 1840 2040
rect 820 1830 880 1840
rect 1340 1830 1400 1840
rect 120 1460 180 1470
rect 60 1260 120 1460
rect 60 1020 180 1260
rect 60 820 120 1020
rect 120 810 180 820
rect 260 1460 320 1470
rect 560 1460 620 1470
rect 1080 1460 1140 1470
rect 1600 1460 1660 1470
rect 320 1260 560 1460
rect 620 1260 1080 1460
rect 1140 1260 1600 1460
rect 260 1020 440 1260
rect 560 1250 620 1260
rect 1080 1250 1140 1260
rect 1600 1250 1660 1260
rect 560 1020 620 1030
rect 1080 1020 1140 1030
rect 1600 1020 1660 1030
rect 320 820 560 1020
rect 620 820 1080 1020
rect 1140 820 1600 1020
rect 260 810 320 820
rect 560 810 620 820
rect 1080 810 1140 820
rect 1600 810 1660 820
rect 820 420 880 430
rect 1340 420 1400 430
rect 1720 420 1920 1840
rect 880 220 1340 420
rect 1400 220 1840 420
rect 820 210 880 220
rect 1340 210 1400 220
rect 1840 210 1920 220
use sky130_fd_pr__pfet_01v8_ACY9XJ#0  sky130_fd_pr__pfet_01v8_ACY9XJ_0
timestamp 1647254192
transform 1 0 216 0 1 1137
box -216 -1137 216 1137
use sky130_fd_pr__pfet_01v8_J24RLQ#0  sky130_fd_pr__pfet_01v8_J24RLQ_0
timestamp 1647254192
transform 1 0 1232 0 1 1137
box -812 -1137 812 1137
<< end >>
