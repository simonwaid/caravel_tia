magic
tech sky130A
magscale 1 2
timestamp 1646921651
<< pwell >>
rect 4410 8570 5630 8630
rect 4410 7700 4470 8570
rect 5570 7700 5630 8570
rect 4410 7550 5630 7700
rect 4410 6680 4470 7550
rect 5570 6680 5630 7550
rect 4410 6620 4550 6680
rect 5500 6620 5630 6680
<< metal1 >>
rect 4504 8630 5390 8632
rect 4410 8570 5630 8630
rect 4410 7700 4470 8570
rect 4504 8566 5390 8570
rect 4590 8340 4600 8510
rect 4660 8340 4670 8510
rect 4790 8340 4800 8510
rect 4860 8340 4870 8510
rect 4980 8340 4990 8510
rect 5050 8340 5060 8510
rect 5170 8340 5180 8510
rect 5240 8340 5250 8510
rect 5360 8340 5370 8510
rect 5430 8340 5440 8510
rect 4500 7740 4510 7910
rect 4570 7740 4580 7910
rect 4690 7740 4700 7910
rect 4760 7740 4770 7910
rect 4880 7740 4890 7910
rect 4950 7740 4960 7910
rect 5070 7740 5080 7910
rect 5140 7740 5150 7910
rect 5270 7740 5280 7910
rect 5340 7740 5350 7910
rect 5460 7740 5470 7910
rect 5530 7740 5540 7910
rect 5570 7700 5630 8570
rect 4410 7550 5630 7700
rect 4410 6680 4470 7550
rect 4590 7330 4600 7500
rect 4660 7330 4670 7500
rect 4790 7330 4800 7500
rect 4860 7330 4870 7500
rect 4980 7330 4990 7500
rect 5050 7330 5060 7500
rect 5170 7330 5180 7500
rect 5240 7330 5250 7500
rect 5360 7330 5370 7500
rect 5430 7330 5440 7500
rect 4500 6730 4510 6900
rect 4570 6730 4580 6900
rect 4690 6730 4700 6900
rect 4760 6730 4770 6900
rect 4880 6730 4890 6900
rect 4950 6730 4960 6900
rect 5070 6730 5080 6900
rect 5140 6730 5150 6900
rect 5270 6730 5280 6900
rect 5340 6730 5350 6900
rect 5460 6730 5470 6900
rect 5530 6730 5540 6900
rect 5570 6680 5630 7550
rect 4410 6620 5630 6680
<< via1 >>
rect 4600 8340 4660 8510
rect 4800 8340 4860 8510
rect 4990 8340 5050 8510
rect 5180 8340 5240 8510
rect 5370 8340 5430 8510
rect 4510 7740 4570 7910
rect 4700 7740 4760 7910
rect 4890 7740 4950 7910
rect 5080 7740 5140 7910
rect 5280 7740 5340 7910
rect 5470 7740 5530 7910
rect 4600 7330 4660 7500
rect 4800 7330 4860 7500
rect 4990 7330 5050 7500
rect 5180 7330 5240 7500
rect 5370 7330 5430 7500
rect 4510 6730 4570 6900
rect 4700 6730 4760 6900
rect 4890 6730 4950 6900
rect 5080 6730 5140 6900
rect 5280 6730 5340 6900
rect 5470 6730 5530 6900
<< metal2 >>
rect 4600 8510 4660 8520
rect 4800 8510 4860 8520
rect 4990 8510 5050 8520
rect 5180 8510 5240 8520
rect 5370 8510 5430 8520
rect 4250 8340 4600 8510
rect 4660 8340 4800 8510
rect 4860 8340 4990 8510
rect 5050 8340 5180 8510
rect 5240 8340 5370 8510
rect 5430 8340 5530 8510
rect 4250 7500 4450 8340
rect 4600 8330 4660 8340
rect 4800 8330 4860 8340
rect 4990 8330 5050 8340
rect 5180 8330 5240 8340
rect 5370 8330 5430 8340
rect 4510 7910 4570 7920
rect 4700 7910 4760 7920
rect 4890 7910 4950 7920
rect 5080 7910 5140 7920
rect 5280 7910 5340 7920
rect 5470 7910 5530 7920
rect 4570 7740 4700 7910
rect 4760 7740 4890 7910
rect 4950 7740 5080 7910
rect 5140 7740 5280 7910
rect 5340 7740 5470 7910
rect 5530 7740 5820 7910
rect 4510 7730 4570 7740
rect 4700 7730 4760 7740
rect 4890 7730 4950 7740
rect 5080 7730 5140 7740
rect 5280 7730 5340 7740
rect 5470 7730 5530 7740
rect 4600 7500 4660 7510
rect 4800 7500 4860 7510
rect 4990 7500 5050 7510
rect 5180 7500 5240 7510
rect 5370 7500 5430 7510
rect 4250 7330 4600 7500
rect 4660 7330 4800 7500
rect 4860 7330 4990 7500
rect 5050 7330 5180 7500
rect 5240 7330 5370 7500
rect 5430 7330 5530 7500
rect 4250 7320 4450 7330
rect 4600 7320 4660 7330
rect 4800 7320 4860 7330
rect 4990 7320 5050 7330
rect 5180 7320 5240 7330
rect 5370 7320 5430 7330
rect 4510 6900 4570 6910
rect 4700 6900 4760 6910
rect 4890 6900 4950 6910
rect 5080 6900 5140 6910
rect 5280 6900 5340 6910
rect 5470 6900 5530 6910
rect 5620 6900 5820 7740
rect 4570 6730 4700 6900
rect 4760 6730 4890 6900
rect 4950 6730 5080 6900
rect 5140 6730 5280 6900
rect 5340 6730 5470 6900
rect 5530 6730 5820 6900
rect 4510 6720 4570 6730
rect 4700 6720 4760 6730
rect 4890 6720 4950 6730
rect 5080 6720 5140 6730
rect 5280 6720 5340 6730
rect 5470 6720 5530 6730
use sky130_fd_pr__nfet_01v8_lvt_26RGPZ  sky130_fd_pr__nfet_01v8_lvt_26RGPZ_0
timestamp 1646921651
transform 1 0 5017 0 1 7629
box -647 -1119 647 1119
<< end >>
