magic
tech sky130A
magscale 1 2
timestamp 1645698808
<< dnwell >>
rect 14640 -8120 18160 -5280
<< nwell >>
rect 14560 -5486 18240 -5200
rect 14560 -7914 14846 -5486
rect 17954 -7914 18240 -5486
rect 14560 -8200 18240 -7914
<< nsubdiff >>
rect 14597 -5257 18203 -5237
rect 14597 -5291 14677 -5257
rect 18123 -5291 18203 -5257
rect 14597 -5311 18203 -5291
rect 14597 -5317 14671 -5311
rect 14597 -8083 14617 -5317
rect 14651 -8083 14671 -5317
rect 14597 -8089 14671 -8083
rect 18129 -5317 18203 -5311
rect 18129 -8083 18149 -5317
rect 18183 -8083 18203 -5317
rect 18129 -8089 18203 -8083
rect 14597 -8109 18203 -8089
rect 14597 -8143 14677 -8109
rect 18123 -8143 18203 -8109
rect 14597 -8163 18203 -8143
<< nsubdiffcont >>
rect 14677 -5291 18123 -5257
rect 14617 -8083 14651 -5317
rect 18149 -8083 18183 -5317
rect 14677 -8143 18123 -8109
<< locali >>
rect 14617 -5291 14677 -5257
rect 18123 -5291 18183 -5257
rect 14617 -5317 14651 -5291
rect 18149 -5317 18183 -5291
rect 14617 -8109 14651 -8083
rect 18149 -8109 18183 -8083
rect 14617 -8143 14677 -8109
rect 18123 -8143 18183 -8109
<< viali >>
rect 18120 -5540 18149 -5340
rect 18149 -5540 18183 -5340
rect 18183 -5540 18200 -5340
rect 14940 -7200 15020 -7000
<< metal1 >>
rect 18114 -5340 18206 -5328
rect 17960 -5540 18120 -5340
rect 18200 -5540 18206 -5340
rect 18114 -5552 18206 -5540
rect 15120 -5740 17700 -5680
rect 15050 -6020 15060 -5820
rect 15140 -6020 15150 -5820
rect 15200 -6640 15280 -5740
rect 15570 -6020 15580 -5820
rect 15660 -6020 15670 -5820
rect 16090 -6020 16100 -5820
rect 16180 -6020 16190 -5820
rect 16610 -6020 16620 -5820
rect 16700 -6020 16710 -5820
rect 17130 -6020 17140 -5820
rect 17220 -6020 17230 -5820
rect 15310 -6580 15320 -6380
rect 15400 -6580 15410 -6380
rect 15830 -6580 15840 -6380
rect 15920 -6580 15930 -6380
rect 16350 -6580 16360 -6380
rect 16440 -6580 16450 -6380
rect 16870 -6580 16880 -6380
rect 16960 -6580 16970 -6380
rect 17370 -6580 17380 -6380
rect 17460 -6580 17470 -6380
rect 17520 -6640 17600 -5740
rect 17650 -6020 17660 -5820
rect 17740 -6020 17750 -5820
rect 14640 -6760 17700 -6640
rect 14934 -7000 15026 -6988
rect 14934 -7020 14940 -7000
rect 14640 -7140 14940 -7020
rect 14934 -7200 14940 -7140
rect 15020 -7200 15026 -7000
rect 14934 -7212 15026 -7200
rect 15050 -7600 15060 -7400
rect 15140 -7600 15150 -7400
rect 15200 -7660 15280 -6760
rect 15310 -7040 15320 -6840
rect 15400 -7040 15410 -6840
rect 15830 -7040 15840 -6840
rect 15920 -7040 15930 -6840
rect 16350 -7040 16360 -6840
rect 16440 -7040 16450 -6840
rect 16870 -7040 16880 -6840
rect 16960 -7040 16970 -6840
rect 17370 -7040 17380 -6840
rect 17460 -7040 17470 -6840
rect 15570 -7600 15580 -7400
rect 15660 -7600 15670 -7400
rect 16090 -7600 16100 -7400
rect 16180 -7600 16190 -7400
rect 16610 -7600 16620 -7400
rect 16700 -7600 16710 -7400
rect 17130 -7600 17140 -7400
rect 17220 -7600 17230 -7400
rect 17520 -7660 17600 -6760
rect 17650 -7600 17660 -7400
rect 17740 -7600 17750 -7400
rect 15120 -7720 17700 -7660
<< via1 >>
rect 15060 -6020 15140 -5820
rect 15580 -6020 15660 -5820
rect 16100 -6020 16180 -5820
rect 16620 -6020 16700 -5820
rect 17140 -6020 17220 -5820
rect 15320 -6580 15400 -6380
rect 15840 -6580 15920 -6380
rect 16360 -6580 16440 -6380
rect 16880 -6580 16960 -6380
rect 17380 -6580 17460 -6380
rect 17660 -6020 17740 -5820
rect 15060 -7600 15140 -7400
rect 15320 -7040 15400 -6840
rect 15840 -7040 15920 -6840
rect 16360 -7040 16440 -6840
rect 16880 -7040 16960 -6840
rect 17380 -7040 17460 -6840
rect 15580 -7600 15660 -7400
rect 16100 -7600 16180 -7400
rect 16620 -7600 16700 -7400
rect 17140 -7600 17220 -7400
rect 17660 -7600 17740 -7400
<< metal2 >>
rect 15060 -5820 15140 -5810
rect 15580 -5820 15660 -5810
rect 16100 -5820 16180 -5810
rect 16620 -5820 16700 -5810
rect 17140 -5820 17220 -5810
rect 17660 -5820 17740 -5810
rect 15140 -6020 15580 -5820
rect 15660 -6020 16100 -5820
rect 16180 -6020 16620 -5820
rect 16700 -6020 17140 -5820
rect 17220 -6020 17660 -5820
rect 15060 -6820 15240 -6020
rect 15580 -6030 15660 -6020
rect 16100 -6030 16180 -6020
rect 16620 -6030 16700 -6020
rect 17140 -6030 17220 -6020
rect 17660 -6030 17740 -6020
rect 14640 -6960 15240 -6820
rect 15060 -7400 15240 -6960
rect 15320 -6380 15400 -6370
rect 15840 -6380 15920 -6370
rect 16360 -6380 16440 -6370
rect 16880 -6380 16960 -6370
rect 17380 -6380 17460 -6370
rect 15400 -6580 15840 -6380
rect 15920 -6580 16360 -6380
rect 16440 -6580 16880 -6380
rect 16960 -6580 17380 -6380
rect 15320 -6600 17460 -6580
rect 15320 -6800 18080 -6600
rect 15320 -6840 17460 -6800
rect 15400 -7040 15840 -6840
rect 15920 -7040 16360 -6840
rect 16440 -7040 16880 -6840
rect 16960 -7040 17380 -6840
rect 15320 -7050 15400 -7040
rect 15840 -7050 15920 -7040
rect 16360 -7050 16440 -7040
rect 16880 -7050 16960 -7040
rect 17380 -7050 17460 -7040
rect 15580 -7400 15660 -7390
rect 16100 -7400 16180 -7390
rect 16620 -7400 16700 -7390
rect 17140 -7400 17220 -7390
rect 17660 -7400 17740 -7390
rect 15140 -7600 15580 -7400
rect 15660 -7600 16100 -7400
rect 16180 -7600 16620 -7400
rect 16700 -7600 17140 -7400
rect 17220 -7600 17660 -7400
rect 15060 -7610 15140 -7600
rect 15580 -7610 15660 -7600
rect 16100 -7610 16180 -7600
rect 16620 -7610 16700 -7600
rect 17140 -7610 17220 -7600
rect 17660 -7610 17740 -7600
use sky130_fd_pr__nfet_01v8_lvt_ZZ3Y87  sky130_fd_pr__nfet_01v8_lvt_ZZ3Y87_0
timestamp 1645633816
transform 1 0 16397 0 1 -6701
box -1457 -1119 1457 1119
<< end >>
