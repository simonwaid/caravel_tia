magic
tech sky130A
timestamp 1647254192
<< nwell >>
rect -1990 -199 1990 199
<< pwell >>
rect -2080 199 2080 289
rect -2080 -199 -1990 199
rect 1990 -199 2080 199
rect -2080 -289 2080 -199
<< mvpsubdiff >>
rect -2062 265 2062 271
rect -2062 248 -2008 265
rect 2008 248 2062 265
rect -2062 242 2062 248
rect -2062 217 -2033 242
rect -2062 -217 -2056 217
rect -2039 -217 -2033 217
rect 2033 217 2062 242
rect -2062 -242 -2033 -217
rect 2033 -217 2039 217
rect 2056 -217 2062 217
rect 2033 -242 2062 -217
rect -2062 -248 2062 -242
rect -2062 -265 -2008 -248
rect 2008 -265 2062 -248
rect -2062 -271 2062 -265
<< mvnsubdiff >>
rect -1957 160 -1625 166
rect -1957 143 -1903 160
rect -1679 143 -1625 160
rect -1957 137 -1625 143
rect -1957 112 -1928 137
rect -1957 -112 -1951 112
rect -1934 -112 -1928 112
rect -1654 112 -1625 137
rect -1957 -137 -1928 -112
rect -1654 -112 -1648 112
rect -1631 -112 -1625 112
rect -1654 -137 -1625 -112
rect -1957 -143 -1625 -137
rect -1957 -160 -1903 -143
rect -1679 -160 -1625 -143
rect -1957 -166 -1625 -160
rect -1559 160 -1227 166
rect -1559 143 -1505 160
rect -1281 143 -1227 160
rect -1559 137 -1227 143
rect -1559 112 -1530 137
rect -1559 -112 -1553 112
rect -1536 -112 -1530 112
rect -1256 112 -1227 137
rect -1559 -137 -1530 -112
rect -1256 -112 -1250 112
rect -1233 -112 -1227 112
rect -1256 -137 -1227 -112
rect -1559 -143 -1227 -137
rect -1559 -160 -1505 -143
rect -1281 -160 -1227 -143
rect -1559 -166 -1227 -160
rect -1161 160 -829 166
rect -1161 143 -1107 160
rect -883 143 -829 160
rect -1161 137 -829 143
rect -1161 112 -1132 137
rect -1161 -112 -1155 112
rect -1138 -112 -1132 112
rect -858 112 -829 137
rect -1161 -137 -1132 -112
rect -858 -112 -852 112
rect -835 -112 -829 112
rect -858 -137 -829 -112
rect -1161 -143 -829 -137
rect -1161 -160 -1107 -143
rect -883 -160 -829 -143
rect -1161 -166 -829 -160
rect -763 160 -431 166
rect -763 143 -709 160
rect -485 143 -431 160
rect -763 137 -431 143
rect -763 112 -734 137
rect -763 -112 -757 112
rect -740 -112 -734 112
rect -460 112 -431 137
rect -763 -137 -734 -112
rect -460 -112 -454 112
rect -437 -112 -431 112
rect -460 -137 -431 -112
rect -763 -143 -431 -137
rect -763 -160 -709 -143
rect -485 -160 -431 -143
rect -763 -166 -431 -160
rect -365 160 -33 166
rect -365 143 -311 160
rect -87 143 -33 160
rect -365 137 -33 143
rect -365 112 -336 137
rect -365 -112 -359 112
rect -342 -112 -336 112
rect -62 112 -33 137
rect -365 -137 -336 -112
rect -62 -112 -56 112
rect -39 -112 -33 112
rect -62 -137 -33 -112
rect -365 -143 -33 -137
rect -365 -160 -311 -143
rect -87 -160 -33 -143
rect -365 -166 -33 -160
rect 33 160 365 166
rect 33 143 87 160
rect 311 143 365 160
rect 33 137 365 143
rect 33 112 62 137
rect 33 -112 39 112
rect 56 -112 62 112
rect 336 112 365 137
rect 33 -137 62 -112
rect 336 -112 342 112
rect 359 -112 365 112
rect 336 -137 365 -112
rect 33 -143 365 -137
rect 33 -160 87 -143
rect 311 -160 365 -143
rect 33 -166 365 -160
rect 431 160 763 166
rect 431 143 485 160
rect 709 143 763 160
rect 431 137 763 143
rect 431 112 460 137
rect 431 -112 437 112
rect 454 -112 460 112
rect 734 112 763 137
rect 431 -137 460 -112
rect 734 -112 740 112
rect 757 -112 763 112
rect 734 -137 763 -112
rect 431 -143 763 -137
rect 431 -160 485 -143
rect 709 -160 763 -143
rect 431 -166 763 -160
rect 829 160 1161 166
rect 829 143 883 160
rect 1107 143 1161 160
rect 829 137 1161 143
rect 829 112 858 137
rect 829 -112 835 112
rect 852 -112 858 112
rect 1132 112 1161 137
rect 829 -137 858 -112
rect 1132 -112 1138 112
rect 1155 -112 1161 112
rect 1132 -137 1161 -112
rect 829 -143 1161 -137
rect 829 -160 883 -143
rect 1107 -160 1161 -143
rect 829 -166 1161 -160
rect 1227 160 1559 166
rect 1227 143 1281 160
rect 1505 143 1559 160
rect 1227 137 1559 143
rect 1227 112 1256 137
rect 1227 -112 1233 112
rect 1250 -112 1256 112
rect 1530 112 1559 137
rect 1227 -137 1256 -112
rect 1530 -112 1536 112
rect 1553 -112 1559 112
rect 1530 -137 1559 -112
rect 1227 -143 1559 -137
rect 1227 -160 1281 -143
rect 1505 -160 1559 -143
rect 1227 -166 1559 -160
rect 1625 160 1957 166
rect 1625 143 1679 160
rect 1903 143 1957 160
rect 1625 137 1957 143
rect 1625 112 1654 137
rect 1625 -112 1631 112
rect 1648 -112 1654 112
rect 1928 112 1957 137
rect 1625 -137 1654 -112
rect 1928 -112 1934 112
rect 1951 -112 1957 112
rect 1928 -137 1957 -112
rect 1625 -143 1957 -137
rect 1625 -160 1679 -143
rect 1903 -160 1957 -143
rect 1625 -166 1957 -160
<< mvpsubdiffcont >>
rect -2008 248 2008 265
rect -2056 -217 -2039 217
rect 2039 -217 2056 217
rect -2008 -265 2008 -248
<< mvnsubdiffcont >>
rect -1903 143 -1679 160
rect -1951 -112 -1934 112
rect -1648 -112 -1631 112
rect -1903 -160 -1679 -143
rect -1505 143 -1281 160
rect -1553 -112 -1536 112
rect -1250 -112 -1233 112
rect -1505 -160 -1281 -143
rect -1107 143 -883 160
rect -1155 -112 -1138 112
rect -852 -112 -835 112
rect -1107 -160 -883 -143
rect -709 143 -485 160
rect -757 -112 -740 112
rect -454 -112 -437 112
rect -709 -160 -485 -143
rect -311 143 -87 160
rect -359 -112 -342 112
rect -56 -112 -39 112
rect -311 -160 -87 -143
rect 87 143 311 160
rect 39 -112 56 112
rect 342 -112 359 112
rect 87 -160 311 -143
rect 485 143 709 160
rect 437 -112 454 112
rect 740 -112 757 112
rect 485 -160 709 -143
rect 883 143 1107 160
rect 835 -112 852 112
rect 1138 -112 1155 112
rect 883 -160 1107 -143
rect 1281 143 1505 160
rect 1233 -112 1250 112
rect 1536 -112 1553 112
rect 1281 -160 1505 -143
rect 1679 143 1903 160
rect 1631 -112 1648 112
rect 1934 -112 1951 112
rect 1679 -160 1903 -143
<< mvpdiode >>
rect -1891 94 -1691 100
rect -1891 -94 -1885 94
rect -1697 -94 -1691 94
rect -1891 -100 -1691 -94
rect -1493 94 -1293 100
rect -1493 -94 -1487 94
rect -1299 -94 -1293 94
rect -1493 -100 -1293 -94
rect -1095 94 -895 100
rect -1095 -94 -1089 94
rect -901 -94 -895 94
rect -1095 -100 -895 -94
rect -697 94 -497 100
rect -697 -94 -691 94
rect -503 -94 -497 94
rect -697 -100 -497 -94
rect -299 94 -99 100
rect -299 -94 -293 94
rect -105 -94 -99 94
rect -299 -100 -99 -94
rect 99 94 299 100
rect 99 -94 105 94
rect 293 -94 299 94
rect 99 -100 299 -94
rect 497 94 697 100
rect 497 -94 503 94
rect 691 -94 697 94
rect 497 -100 697 -94
rect 895 94 1095 100
rect 895 -94 901 94
rect 1089 -94 1095 94
rect 895 -100 1095 -94
rect 1293 94 1493 100
rect 1293 -94 1299 94
rect 1487 -94 1493 94
rect 1293 -100 1493 -94
rect 1691 94 1891 100
rect 1691 -94 1697 94
rect 1885 -94 1891 94
rect 1691 -100 1891 -94
<< mvpdiodec >>
rect -1885 -94 -1697 94
rect -1487 -94 -1299 94
rect -1089 -94 -901 94
rect -691 -94 -503 94
rect -293 -94 -105 94
rect 105 -94 293 94
rect 503 -94 691 94
rect 901 -94 1089 94
rect 1299 -94 1487 94
rect 1697 -94 1885 94
<< locali >>
rect -2056 248 -2008 265
rect 2008 248 2056 265
rect -2056 217 -2039 248
rect 2039 217 2056 248
rect -1951 143 -1903 160
rect -1679 143 -1631 160
rect -1951 112 -1934 143
rect -1648 112 -1631 143
rect -1893 -94 -1885 94
rect -1697 -94 -1689 94
rect -1951 -143 -1934 -112
rect -1648 -143 -1631 -112
rect -1951 -160 -1903 -143
rect -1679 -160 -1631 -143
rect -1553 143 -1505 160
rect -1281 143 -1233 160
rect -1553 112 -1536 143
rect -1250 112 -1233 143
rect -1495 -94 -1487 94
rect -1299 -94 -1291 94
rect -1553 -143 -1536 -112
rect -1250 -143 -1233 -112
rect -1553 -160 -1505 -143
rect -1281 -160 -1233 -143
rect -1155 143 -1107 160
rect -883 143 -835 160
rect -1155 112 -1138 143
rect -852 112 -835 143
rect -1097 -94 -1089 94
rect -901 -94 -893 94
rect -1155 -143 -1138 -112
rect -852 -143 -835 -112
rect -1155 -160 -1107 -143
rect -883 -160 -835 -143
rect -757 143 -709 160
rect -485 143 -437 160
rect -757 112 -740 143
rect -454 112 -437 143
rect -699 -94 -691 94
rect -503 -94 -495 94
rect -757 -143 -740 -112
rect -454 -143 -437 -112
rect -757 -160 -709 -143
rect -485 -160 -437 -143
rect -359 143 -311 160
rect -87 143 -39 160
rect -359 112 -342 143
rect -56 112 -39 143
rect -301 -94 -293 94
rect -105 -94 -97 94
rect -359 -143 -342 -112
rect -56 -143 -39 -112
rect -359 -160 -311 -143
rect -87 -160 -39 -143
rect 39 143 87 160
rect 311 143 359 160
rect 39 112 56 143
rect 342 112 359 143
rect 97 -94 105 94
rect 293 -94 301 94
rect 39 -143 56 -112
rect 342 -143 359 -112
rect 39 -160 87 -143
rect 311 -160 359 -143
rect 437 143 485 160
rect 709 143 757 160
rect 437 112 454 143
rect 740 112 757 143
rect 495 -94 503 94
rect 691 -94 699 94
rect 437 -143 454 -112
rect 740 -143 757 -112
rect 437 -160 485 -143
rect 709 -160 757 -143
rect 835 143 883 160
rect 1107 143 1155 160
rect 835 112 852 143
rect 1138 112 1155 143
rect 893 -94 901 94
rect 1089 -94 1097 94
rect 835 -143 852 -112
rect 1138 -143 1155 -112
rect 835 -160 883 -143
rect 1107 -160 1155 -143
rect 1233 143 1281 160
rect 1505 143 1553 160
rect 1233 112 1250 143
rect 1536 112 1553 143
rect 1291 -94 1299 94
rect 1487 -94 1495 94
rect 1233 -143 1250 -112
rect 1536 -143 1553 -112
rect 1233 -160 1281 -143
rect 1505 -160 1553 -143
rect 1631 143 1679 160
rect 1903 143 1951 160
rect 1631 112 1648 143
rect 1934 112 1951 143
rect 1689 -94 1697 94
rect 1885 -94 1893 94
rect 1631 -143 1648 -112
rect 1934 -143 1951 -112
rect 1631 -160 1679 -143
rect 1903 -160 1951 -143
rect -2056 -248 -2039 -217
rect 2039 -248 2056 -217
rect -2056 -265 -2008 -248
rect 2008 -265 2056 -248
<< viali >>
rect -1885 -94 -1697 94
rect -1487 -94 -1299 94
rect -1089 -94 -901 94
rect -691 -94 -503 94
rect -293 -94 -105 94
rect 105 -94 293 94
rect 503 -94 691 94
rect 901 -94 1089 94
rect 1299 -94 1487 94
rect 1697 -94 1885 94
<< metal1 >>
rect -1891 94 -1691 97
rect -1891 -94 -1885 94
rect -1697 -94 -1691 94
rect -1891 -97 -1691 -94
rect -1493 94 -1293 97
rect -1493 -94 -1487 94
rect -1299 -94 -1293 94
rect -1493 -97 -1293 -94
rect -1095 94 -895 97
rect -1095 -94 -1089 94
rect -901 -94 -895 94
rect -1095 -97 -895 -94
rect -697 94 -497 97
rect -697 -94 -691 94
rect -503 -94 -497 94
rect -697 -97 -497 -94
rect -299 94 -99 97
rect -299 -94 -293 94
rect -105 -94 -99 94
rect -299 -97 -99 -94
rect 99 94 299 97
rect 99 -94 105 94
rect 293 -94 299 94
rect 99 -97 299 -94
rect 497 94 697 97
rect 497 -94 503 94
rect 691 -94 697 94
rect 497 -97 697 -94
rect 895 94 1095 97
rect 895 -94 901 94
rect 1089 -94 1095 94
rect 895 -97 1095 -94
rect 1293 94 1493 97
rect 1293 -94 1299 94
rect 1487 -94 1493 94
rect 1293 -97 1493 -94
rect 1691 94 1891 97
rect 1691 -94 1697 94
rect 1885 -94 1891 94
rect 1691 -97 1891 -94
<< properties >>
string FIXED_BBOX 1639 -151 1942 151
string gencell sky130_fd_pr__diode_pd2nw_11v0
string library sky130
string parameters w 2 l 2 area 4.0 peri 8.0 nx 10 ny 1 dummy 0 lmin 0.45 wmin 0.45 elc 1 erc 1 etc 1 ebc 1 glc 1 grc 1 gtc 1 gbc 1 doverlap 0 compatible {sky130_fd_pr__diode_pd2nw_05v5 sky130_fd_pr__diode_pd2nw_05v5_lvt  sky130_fd_pr__diode_pd2nw_05v5_hvt sky130_fd_pr__diode_pd2nw_11v0} full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
