magic
tech sky130A
magscale 1 2
timestamp 1647255486
<< dnwell >>
rect 2094 -710 4374 1210
rect 2094 -7780 4374 -5860
<< nwell >>
rect -1326 2112 2276 2764
rect -1326 1290 4188 2112
rect 2014 1004 4454 1290
rect 2014 -504 2300 1004
rect 4168 -504 4454 1004
rect 2014 -790 4454 -504
rect -1326 -4958 2276 -4306
rect -1326 -5780 4188 -4958
rect 2014 -6066 4454 -5780
rect 2014 -7574 2300 -6066
rect 4168 -7574 4454 -6066
rect 2014 -7860 4454 -7574
rect 1560 -11040 2226 -9804
rect 2480 -11040 3146 -9804
rect 3400 -11040 4066 -9804
rect 4320 -11040 4986 -9804
rect 5240 -11040 5906 -9804
rect 6180 -10530 6772 -9992
<< pwell >>
rect -1326 1220 1458 1288
rect -1326 1140 1464 1220
rect -1326 640 1458 1140
rect -1336 490 1464 640
rect -1326 30 1458 490
rect -1336 -30 1464 30
rect -1326 -150 1458 -30
rect -1326 -260 1458 -156
rect -1336 -270 1458 -260
rect -1336 -330 1464 -270
rect -1326 -800 1458 -330
rect 2334 -470 4138 968
rect -1336 -810 1464 -800
rect -1336 -950 2950 -810
rect -1326 -1576 1458 -950
rect -1346 -1594 1458 -1576
rect -1346 -4250 1388 -1594
rect 1464 -1630 2950 -950
rect 1464 -2450 3346 -1630
rect -1326 -5850 1458 -5782
rect -1326 -5930 1464 -5850
rect -1326 -6430 1458 -5930
rect -1336 -6580 1464 -6430
rect -1326 -7040 1458 -6580
rect -1336 -7100 1464 -7040
rect -1326 -7220 1458 -7100
rect -1326 -7330 1458 -7226
rect -1336 -7340 1458 -7330
rect -1336 -7400 1464 -7340
rect -1326 -7870 1458 -7400
rect 2334 -7540 4138 -6102
rect -1336 -7880 1464 -7870
rect -1336 -8020 2950 -7880
rect -1326 -8646 1458 -8020
rect -1346 -8664 1458 -8646
rect -1346 -11320 1388 -8664
rect 1464 -8700 2950 -8020
rect 3360 -8700 4846 -7880
rect 1464 -9520 3346 -8700
rect 3360 -9520 5242 -8700
rect 5310 -9520 6124 -8700
rect 1450 -9804 6016 -9694
rect 1450 -11040 1560 -9804
rect 2226 -11040 2480 -9804
rect 3146 -11040 3400 -9804
rect 4066 -11040 4320 -9804
rect 4986 -11040 5240 -9804
rect 5906 -11040 6016 -9804
rect 1450 -11150 6016 -11040
rect 6180 -11080 6772 -10560
<< nmos >>
rect 1664 -1420 1694 -1020
rect 1760 -1420 1790 -1020
rect 1856 -1420 1886 -1020
rect 1952 -1420 1982 -1020
rect 2048 -1420 2078 -1020
rect 2144 -1420 2174 -1020
rect 2240 -1420 2270 -1020
rect 2336 -1420 2366 -1020
rect 2432 -1420 2462 -1020
rect 2528 -1420 2558 -1020
rect 2624 -1420 2654 -1020
rect 2720 -1420 2750 -1020
rect -1146 -2186 -1116 -1786
rect -1050 -2186 -1020 -1786
rect -954 -2186 -924 -1786
rect -858 -2186 -828 -1786
rect -762 -2186 -732 -1786
rect -666 -2186 -636 -1786
rect -570 -2186 -540 -1786
rect -474 -2186 -444 -1786
rect -378 -2186 -348 -1786
rect -282 -2186 -252 -1786
rect -186 -2186 -156 -1786
rect -90 -2186 -60 -1786
rect 6 -2186 36 -1786
rect 102 -2186 132 -1786
rect 198 -2186 228 -1786
rect 294 -2186 324 -1786
rect 390 -2186 420 -1786
rect 486 -2186 516 -1786
rect 582 -2186 612 -1786
rect 678 -2186 708 -1786
rect 774 -2186 804 -1786
rect 870 -2186 900 -1786
rect 966 -2186 996 -1786
rect 1062 -2186 1092 -1786
rect 1158 -2186 1188 -1786
rect -1146 -2804 -1116 -2404
rect -1050 -2804 -1020 -2404
rect -954 -2804 -924 -2404
rect -858 -2804 -828 -2404
rect -762 -2804 -732 -2404
rect -666 -2804 -636 -2404
rect -570 -2804 -540 -2404
rect -474 -2804 -444 -2404
rect -378 -2804 -348 -2404
rect -282 -2804 -252 -2404
rect -186 -2804 -156 -2404
rect -90 -2804 -60 -2404
rect 6 -2804 36 -2404
rect 102 -2804 132 -2404
rect 198 -2804 228 -2404
rect 294 -2804 324 -2404
rect 390 -2804 420 -2404
rect 486 -2804 516 -2404
rect 582 -2804 612 -2404
rect 678 -2804 708 -2404
rect 774 -2804 804 -2404
rect 870 -2804 900 -2404
rect 966 -2804 996 -2404
rect 1062 -2804 1092 -2404
rect 1158 -2804 1188 -2404
rect -1146 -3422 -1116 -3022
rect -1050 -3422 -1020 -3022
rect -954 -3422 -924 -3022
rect -858 -3422 -828 -3022
rect -762 -3422 -732 -3022
rect -666 -3422 -636 -3022
rect -570 -3422 -540 -3022
rect -474 -3422 -444 -3022
rect -378 -3422 -348 -3022
rect -282 -3422 -252 -3022
rect -186 -3422 -156 -3022
rect -90 -3422 -60 -3022
rect 6 -3422 36 -3022
rect 102 -3422 132 -3022
rect 198 -3422 228 -3022
rect 294 -3422 324 -3022
rect 390 -3422 420 -3022
rect 486 -3422 516 -3022
rect 582 -3422 612 -3022
rect 678 -3422 708 -3022
rect 774 -3422 804 -3022
rect 870 -3422 900 -3022
rect 966 -3422 996 -3022
rect 1062 -3422 1092 -3022
rect 1158 -3422 1188 -3022
rect -1146 -4040 -1116 -3640
rect -1050 -4040 -1020 -3640
rect -954 -4040 -924 -3640
rect -858 -4040 -828 -3640
rect -762 -4040 -732 -3640
rect -666 -4040 -636 -3640
rect -570 -4040 -540 -3640
rect -474 -4040 -444 -3640
rect -378 -4040 -348 -3640
rect -282 -4040 -252 -3640
rect -186 -4040 -156 -3640
rect -90 -4040 -60 -3640
rect 6 -4040 36 -3640
rect 102 -4040 132 -3640
rect 198 -4040 228 -3640
rect 294 -4040 324 -3640
rect 390 -4040 420 -3640
rect 486 -4040 516 -3640
rect 582 -4040 612 -3640
rect 678 -4040 708 -3640
rect 774 -4040 804 -3640
rect 870 -4040 900 -3640
rect 966 -4040 996 -3640
rect 1062 -4040 1092 -3640
rect 1158 -4040 1188 -3640
rect 1660 -2240 1860 -1840
rect 1918 -2240 2118 -1840
rect 2176 -2240 2376 -1840
rect 2434 -2240 2634 -1840
rect 2692 -2240 2892 -1840
rect 2950 -2240 3150 -1840
rect 1664 -8490 1694 -8090
rect 1760 -8490 1790 -8090
rect 1856 -8490 1886 -8090
rect 1952 -8490 1982 -8090
rect 2048 -8490 2078 -8090
rect 2144 -8490 2174 -8090
rect 2240 -8490 2270 -8090
rect 2336 -8490 2366 -8090
rect 2432 -8490 2462 -8090
rect 2528 -8490 2558 -8090
rect 2624 -8490 2654 -8090
rect 2720 -8490 2750 -8090
rect 3560 -8490 3590 -8090
rect 3656 -8490 3686 -8090
rect 3752 -8490 3782 -8090
rect 3848 -8490 3878 -8090
rect 3944 -8490 3974 -8090
rect 4040 -8490 4070 -8090
rect 4136 -8490 4166 -8090
rect 4232 -8490 4262 -8090
rect 4328 -8490 4358 -8090
rect 4424 -8490 4454 -8090
rect 4520 -8490 4550 -8090
rect 4616 -8490 4646 -8090
rect -1146 -9256 -1116 -8856
rect -1050 -9256 -1020 -8856
rect -954 -9256 -924 -8856
rect -858 -9256 -828 -8856
rect -762 -9256 -732 -8856
rect -666 -9256 -636 -8856
rect -570 -9256 -540 -8856
rect -474 -9256 -444 -8856
rect -378 -9256 -348 -8856
rect -282 -9256 -252 -8856
rect -186 -9256 -156 -8856
rect -90 -9256 -60 -8856
rect 6 -9256 36 -8856
rect 102 -9256 132 -8856
rect 198 -9256 228 -8856
rect 294 -9256 324 -8856
rect 390 -9256 420 -8856
rect 486 -9256 516 -8856
rect 582 -9256 612 -8856
rect 678 -9256 708 -8856
rect 774 -9256 804 -8856
rect 870 -9256 900 -8856
rect 966 -9256 996 -8856
rect 1062 -9256 1092 -8856
rect 1158 -9256 1188 -8856
rect -1146 -9874 -1116 -9474
rect -1050 -9874 -1020 -9474
rect -954 -9874 -924 -9474
rect -858 -9874 -828 -9474
rect -762 -9874 -732 -9474
rect -666 -9874 -636 -9474
rect -570 -9874 -540 -9474
rect -474 -9874 -444 -9474
rect -378 -9874 -348 -9474
rect -282 -9874 -252 -9474
rect -186 -9874 -156 -9474
rect -90 -9874 -60 -9474
rect 6 -9874 36 -9474
rect 102 -9874 132 -9474
rect 198 -9874 228 -9474
rect 294 -9874 324 -9474
rect 390 -9874 420 -9474
rect 486 -9874 516 -9474
rect 582 -9874 612 -9474
rect 678 -9874 708 -9474
rect 774 -9874 804 -9474
rect 870 -9874 900 -9474
rect 966 -9874 996 -9474
rect 1062 -9874 1092 -9474
rect 1158 -9874 1188 -9474
rect -1146 -10492 -1116 -10092
rect -1050 -10492 -1020 -10092
rect -954 -10492 -924 -10092
rect -858 -10492 -828 -10092
rect -762 -10492 -732 -10092
rect -666 -10492 -636 -10092
rect -570 -10492 -540 -10092
rect -474 -10492 -444 -10092
rect -378 -10492 -348 -10092
rect -282 -10492 -252 -10092
rect -186 -10492 -156 -10092
rect -90 -10492 -60 -10092
rect 6 -10492 36 -10092
rect 102 -10492 132 -10092
rect 198 -10492 228 -10092
rect 294 -10492 324 -10092
rect 390 -10492 420 -10092
rect 486 -10492 516 -10092
rect 582 -10492 612 -10092
rect 678 -10492 708 -10092
rect 774 -10492 804 -10092
rect 870 -10492 900 -10092
rect 966 -10492 996 -10092
rect 1062 -10492 1092 -10092
rect 1158 -10492 1188 -10092
rect -1146 -11110 -1116 -10710
rect -1050 -11110 -1020 -10710
rect -954 -11110 -924 -10710
rect -858 -11110 -828 -10710
rect -762 -11110 -732 -10710
rect -666 -11110 -636 -10710
rect -570 -11110 -540 -10710
rect -474 -11110 -444 -10710
rect -378 -11110 -348 -10710
rect -282 -11110 -252 -10710
rect -186 -11110 -156 -10710
rect -90 -11110 -60 -10710
rect 6 -11110 36 -10710
rect 102 -11110 132 -10710
rect 198 -11110 228 -10710
rect 294 -11110 324 -10710
rect 390 -11110 420 -10710
rect 486 -11110 516 -10710
rect 582 -11110 612 -10710
rect 678 -11110 708 -10710
rect 774 -11110 804 -10710
rect 870 -11110 900 -10710
rect 966 -11110 996 -10710
rect 1062 -11110 1092 -10710
rect 1158 -11110 1188 -10710
rect 1660 -9310 1860 -8910
rect 1918 -9310 2118 -8910
rect 2176 -9310 2376 -8910
rect 2434 -9310 2634 -8910
rect 2692 -9310 2892 -8910
rect 2950 -9310 3150 -8910
rect 3556 -9310 3756 -8910
rect 3814 -9310 4014 -8910
rect 4072 -9310 4272 -8910
rect 4330 -9310 4530 -8910
rect 4588 -9310 4788 -8910
rect 4846 -9310 5046 -8910
rect 5510 -9310 5540 -8910
rect 5606 -9310 5636 -8910
rect 5702 -9310 5732 -8910
rect 5798 -9310 5828 -8910
rect 5894 -9310 5924 -8910
rect 6376 -10870 6576 -10770
<< pmos >>
rect -1130 2145 -1090 2545
rect -1032 2145 -992 2545
rect -934 2145 -894 2545
rect -836 2145 -796 2545
rect -738 2145 -698 2545
rect -640 2145 -600 2545
rect -542 2145 -502 2545
rect -444 2145 -404 2545
rect -346 2145 -306 2545
rect -248 2145 -208 2545
rect -150 2145 -110 2545
rect -52 2145 -12 2545
rect 46 2145 86 2545
rect 144 2145 184 2545
rect 242 2145 282 2545
rect -1130 1509 -1090 1909
rect -1032 1509 -992 1909
rect -934 1509 -894 1909
rect -836 1509 -796 1909
rect -738 1509 -698 1909
rect -640 1509 -600 1909
rect -542 1509 -502 1909
rect -444 1509 -404 1909
rect -346 1509 -306 1909
rect -248 1509 -208 1909
rect -150 1509 -110 1909
rect -52 1509 -12 1909
rect 46 1509 86 1909
rect 144 1509 184 1909
rect 242 1509 282 1909
rect 668 2145 708 2545
rect 766 2145 806 2545
rect 864 2145 904 2545
rect 962 2145 1002 2545
rect 1060 2145 1100 2545
rect 1158 2145 1198 2545
rect 1256 2145 1296 2545
rect 1354 2145 1394 2545
rect 1452 2145 1492 2545
rect 1550 2145 1590 2545
rect 1648 2145 1688 2545
rect 1746 2145 1786 2545
rect 1844 2145 1884 2545
rect 1942 2145 1982 2545
rect 2040 2145 2080 2545
rect 668 1509 708 1909
rect 766 1509 806 1909
rect 864 1509 904 1909
rect 962 1509 1002 1909
rect 1060 1509 1100 1909
rect 1158 1509 1198 1909
rect 1256 1509 1296 1909
rect 1354 1509 1394 1909
rect 1452 1509 1492 1909
rect 1550 1509 1590 1909
rect 1648 1509 1688 1909
rect 1746 1509 1786 1909
rect 1844 1509 1884 1909
rect 1942 1509 1982 1909
rect 2040 1509 2080 1909
rect 2470 1493 2570 1893
rect 2628 1493 2728 1893
rect 2786 1493 2886 1893
rect 2944 1493 3044 1893
rect 3102 1493 3202 1893
rect 3260 1493 3360 1893
rect 3418 1493 3518 1893
rect 3576 1493 3676 1893
rect 3734 1493 3834 1893
rect 3892 1493 3992 1893
rect -1130 -4925 -1090 -4525
rect -1032 -4925 -992 -4525
rect -934 -4925 -894 -4525
rect -836 -4925 -796 -4525
rect -738 -4925 -698 -4525
rect -640 -4925 -600 -4525
rect -542 -4925 -502 -4525
rect -444 -4925 -404 -4525
rect -346 -4925 -306 -4525
rect -248 -4925 -208 -4525
rect -150 -4925 -110 -4525
rect -52 -4925 -12 -4525
rect 46 -4925 86 -4525
rect 144 -4925 184 -4525
rect 242 -4925 282 -4525
rect -1130 -5561 -1090 -5161
rect -1032 -5561 -992 -5161
rect -934 -5561 -894 -5161
rect -836 -5561 -796 -5161
rect -738 -5561 -698 -5161
rect -640 -5561 -600 -5161
rect -542 -5561 -502 -5161
rect -444 -5561 -404 -5161
rect -346 -5561 -306 -5161
rect -248 -5561 -208 -5161
rect -150 -5561 -110 -5161
rect -52 -5561 -12 -5161
rect 46 -5561 86 -5161
rect 144 -5561 184 -5161
rect 242 -5561 282 -5161
rect 668 -4925 708 -4525
rect 766 -4925 806 -4525
rect 864 -4925 904 -4525
rect 962 -4925 1002 -4525
rect 1060 -4925 1100 -4525
rect 1158 -4925 1198 -4525
rect 1256 -4925 1296 -4525
rect 1354 -4925 1394 -4525
rect 1452 -4925 1492 -4525
rect 1550 -4925 1590 -4525
rect 1648 -4925 1688 -4525
rect 1746 -4925 1786 -4525
rect 1844 -4925 1884 -4525
rect 1942 -4925 1982 -4525
rect 2040 -4925 2080 -4525
rect 668 -5561 708 -5161
rect 766 -5561 806 -5161
rect 864 -5561 904 -5161
rect 962 -5561 1002 -5161
rect 1060 -5561 1100 -5161
rect 1158 -5561 1198 -5161
rect 1256 -5561 1296 -5161
rect 1354 -5561 1394 -5161
rect 1452 -5561 1492 -5161
rect 1550 -5561 1590 -5161
rect 1648 -5561 1688 -5161
rect 1746 -5561 1786 -5161
rect 1844 -5561 1884 -5161
rect 1942 -5561 1982 -5161
rect 2040 -5561 2080 -5161
rect 2470 -5577 2570 -5177
rect 2628 -5577 2728 -5177
rect 2786 -5577 2886 -5177
rect 2944 -5577 3044 -5177
rect 3102 -5577 3202 -5177
rect 3260 -5577 3360 -5177
rect 3418 -5577 3518 -5177
rect 3576 -5577 3676 -5177
rect 3734 -5577 3834 -5177
rect 3892 -5577 3992 -5177
rect 6376 -10311 6576 -10211
<< varactor >>
rect 1693 -10922 2093 -9922
rect 2613 -10922 3013 -9922
rect 3533 -10922 3933 -9922
rect 4453 -10922 4853 -9922
rect 5373 -10922 5773 -9922
<< nmoslvt >>
rect -1130 678 -1090 1078
rect -1032 678 -992 1078
rect -934 678 -894 1078
rect -836 678 -796 1078
rect -738 678 -698 1078
rect -640 678 -600 1078
rect -542 678 -502 1078
rect -444 678 -404 1078
rect -346 678 -306 1078
rect -248 678 -208 1078
rect -150 678 -110 1078
rect -52 678 -12 1078
rect 46 678 86 1078
rect 144 678 184 1078
rect 242 678 282 1078
rect 340 678 380 1078
rect 438 678 478 1078
rect 536 678 576 1078
rect 634 678 674 1078
rect 732 678 772 1078
rect 830 678 870 1078
rect 928 678 968 1078
rect 1026 678 1066 1078
rect 1124 678 1164 1078
rect 1222 678 1262 1078
rect -1130 60 -1090 460
rect -1032 60 -992 460
rect -934 60 -894 460
rect -836 60 -796 460
rect -738 60 -698 460
rect -640 60 -600 460
rect -542 60 -502 460
rect -444 60 -404 460
rect -346 60 -306 460
rect -248 60 -208 460
rect -150 60 -110 460
rect -52 60 -12 460
rect 46 60 86 460
rect 144 60 184 460
rect 242 60 282 460
rect 340 60 380 460
rect 438 60 478 460
rect 536 60 576 460
rect 634 60 674 460
rect 732 60 772 460
rect 830 60 870 460
rect 928 60 968 460
rect 1026 60 1066 460
rect 1124 60 1164 460
rect 1222 60 1262 460
rect -1130 -766 -1090 -366
rect -1032 -766 -992 -366
rect -934 -766 -894 -366
rect -836 -766 -796 -366
rect -738 -766 -698 -366
rect -640 -766 -600 -366
rect -542 -766 -502 -366
rect -444 -766 -404 -366
rect -346 -766 -306 -366
rect -248 -766 -208 -366
rect -150 -766 -110 -366
rect -52 -766 -12 -366
rect 46 -766 86 -366
rect 144 -766 184 -366
rect 242 -766 282 -366
rect 340 -766 380 -366
rect 438 -766 478 -366
rect 536 -766 576 -366
rect 634 -766 674 -366
rect 732 -766 772 -366
rect 830 -766 870 -366
rect 928 -766 968 -366
rect 1026 -766 1066 -366
rect 1124 -766 1164 -366
rect 1222 -766 1262 -366
rect -1130 -1384 -1090 -984
rect -1032 -1384 -992 -984
rect -934 -1384 -894 -984
rect -836 -1384 -796 -984
rect -738 -1384 -698 -984
rect -640 -1384 -600 -984
rect -542 -1384 -502 -984
rect -444 -1384 -404 -984
rect -346 -1384 -306 -984
rect -248 -1384 -208 -984
rect -150 -1384 -110 -984
rect -52 -1384 -12 -984
rect 46 -1384 86 -984
rect 144 -1384 184 -984
rect 242 -1384 282 -984
rect 340 -1384 380 -984
rect 438 -1384 478 -984
rect 536 -1384 576 -984
rect 634 -1384 674 -984
rect 732 -1384 772 -984
rect 830 -1384 870 -984
rect 928 -1384 968 -984
rect 1026 -1384 1066 -984
rect 1124 -1384 1164 -984
rect 1222 -1384 1262 -984
rect 2530 358 2570 758
rect 2628 358 2668 758
rect 2726 358 2766 758
rect 2824 358 2864 758
rect 2922 358 2962 758
rect 3020 358 3060 758
rect 3118 358 3158 758
rect 3216 358 3256 758
rect 3314 358 3354 758
rect 3412 358 3452 758
rect 3510 358 3550 758
rect 3608 358 3648 758
rect 3706 358 3746 758
rect 3804 358 3844 758
rect 3902 358 3942 758
rect 2530 -260 2570 140
rect 2628 -260 2668 140
rect 2726 -260 2766 140
rect 2824 -260 2864 140
rect 2922 -260 2962 140
rect 3020 -260 3060 140
rect 3118 -260 3158 140
rect 3216 -260 3256 140
rect 3314 -260 3354 140
rect 3412 -260 3452 140
rect 3510 -260 3550 140
rect 3608 -260 3648 140
rect 3706 -260 3746 140
rect 3804 -260 3844 140
rect 3902 -260 3942 140
rect -1130 -6392 -1090 -5992
rect -1032 -6392 -992 -5992
rect -934 -6392 -894 -5992
rect -836 -6392 -796 -5992
rect -738 -6392 -698 -5992
rect -640 -6392 -600 -5992
rect -542 -6392 -502 -5992
rect -444 -6392 -404 -5992
rect -346 -6392 -306 -5992
rect -248 -6392 -208 -5992
rect -150 -6392 -110 -5992
rect -52 -6392 -12 -5992
rect 46 -6392 86 -5992
rect 144 -6392 184 -5992
rect 242 -6392 282 -5992
rect 340 -6392 380 -5992
rect 438 -6392 478 -5992
rect 536 -6392 576 -5992
rect 634 -6392 674 -5992
rect 732 -6392 772 -5992
rect 830 -6392 870 -5992
rect 928 -6392 968 -5992
rect 1026 -6392 1066 -5992
rect 1124 -6392 1164 -5992
rect 1222 -6392 1262 -5992
rect -1130 -7010 -1090 -6610
rect -1032 -7010 -992 -6610
rect -934 -7010 -894 -6610
rect -836 -7010 -796 -6610
rect -738 -7010 -698 -6610
rect -640 -7010 -600 -6610
rect -542 -7010 -502 -6610
rect -444 -7010 -404 -6610
rect -346 -7010 -306 -6610
rect -248 -7010 -208 -6610
rect -150 -7010 -110 -6610
rect -52 -7010 -12 -6610
rect 46 -7010 86 -6610
rect 144 -7010 184 -6610
rect 242 -7010 282 -6610
rect 340 -7010 380 -6610
rect 438 -7010 478 -6610
rect 536 -7010 576 -6610
rect 634 -7010 674 -6610
rect 732 -7010 772 -6610
rect 830 -7010 870 -6610
rect 928 -7010 968 -6610
rect 1026 -7010 1066 -6610
rect 1124 -7010 1164 -6610
rect 1222 -7010 1262 -6610
rect -1130 -7836 -1090 -7436
rect -1032 -7836 -992 -7436
rect -934 -7836 -894 -7436
rect -836 -7836 -796 -7436
rect -738 -7836 -698 -7436
rect -640 -7836 -600 -7436
rect -542 -7836 -502 -7436
rect -444 -7836 -404 -7436
rect -346 -7836 -306 -7436
rect -248 -7836 -208 -7436
rect -150 -7836 -110 -7436
rect -52 -7836 -12 -7436
rect 46 -7836 86 -7436
rect 144 -7836 184 -7436
rect 242 -7836 282 -7436
rect 340 -7836 380 -7436
rect 438 -7836 478 -7436
rect 536 -7836 576 -7436
rect 634 -7836 674 -7436
rect 732 -7836 772 -7436
rect 830 -7836 870 -7436
rect 928 -7836 968 -7436
rect 1026 -7836 1066 -7436
rect 1124 -7836 1164 -7436
rect 1222 -7836 1262 -7436
rect -1130 -8454 -1090 -8054
rect -1032 -8454 -992 -8054
rect -934 -8454 -894 -8054
rect -836 -8454 -796 -8054
rect -738 -8454 -698 -8054
rect -640 -8454 -600 -8054
rect -542 -8454 -502 -8054
rect -444 -8454 -404 -8054
rect -346 -8454 -306 -8054
rect -248 -8454 -208 -8054
rect -150 -8454 -110 -8054
rect -52 -8454 -12 -8054
rect 46 -8454 86 -8054
rect 144 -8454 184 -8054
rect 242 -8454 282 -8054
rect 340 -8454 380 -8054
rect 438 -8454 478 -8054
rect 536 -8454 576 -8054
rect 634 -8454 674 -8054
rect 732 -8454 772 -8054
rect 830 -8454 870 -8054
rect 928 -8454 968 -8054
rect 1026 -8454 1066 -8054
rect 1124 -8454 1164 -8054
rect 1222 -8454 1262 -8054
rect 2530 -6712 2570 -6312
rect 2628 -6712 2668 -6312
rect 2726 -6712 2766 -6312
rect 2824 -6712 2864 -6312
rect 2922 -6712 2962 -6312
rect 3020 -6712 3060 -6312
rect 3118 -6712 3158 -6312
rect 3216 -6712 3256 -6312
rect 3314 -6712 3354 -6312
rect 3412 -6712 3452 -6312
rect 3510 -6712 3550 -6312
rect 3608 -6712 3648 -6312
rect 3706 -6712 3746 -6312
rect 3804 -6712 3844 -6312
rect 3902 -6712 3942 -6312
rect 2530 -7330 2570 -6930
rect 2628 -7330 2668 -6930
rect 2726 -7330 2766 -6930
rect 2824 -7330 2864 -6930
rect 2922 -7330 2962 -6930
rect 3020 -7330 3060 -6930
rect 3118 -7330 3158 -6930
rect 3216 -7330 3256 -6930
rect 3314 -7330 3354 -6930
rect 3412 -7330 3452 -6930
rect 3510 -7330 3550 -6930
rect 3608 -7330 3648 -6930
rect 3706 -7330 3746 -6930
rect 3804 -7330 3844 -6930
rect 3902 -7330 3942 -6930
<< ndiff >>
rect -1188 1066 -1130 1078
rect -1188 690 -1176 1066
rect -1142 690 -1130 1066
rect -1188 678 -1130 690
rect -1090 1066 -1032 1078
rect -1090 690 -1078 1066
rect -1044 690 -1032 1066
rect -1090 678 -1032 690
rect -992 1066 -934 1078
rect -992 690 -980 1066
rect -946 690 -934 1066
rect -992 678 -934 690
rect -894 1066 -836 1078
rect -894 690 -882 1066
rect -848 690 -836 1066
rect -894 678 -836 690
rect -796 1066 -738 1078
rect -796 690 -784 1066
rect -750 690 -738 1066
rect -796 678 -738 690
rect -698 1066 -640 1078
rect -698 690 -686 1066
rect -652 690 -640 1066
rect -698 678 -640 690
rect -600 1066 -542 1078
rect -600 690 -588 1066
rect -554 690 -542 1066
rect -600 678 -542 690
rect -502 1066 -444 1078
rect -502 690 -490 1066
rect -456 690 -444 1066
rect -502 678 -444 690
rect -404 1066 -346 1078
rect -404 690 -392 1066
rect -358 690 -346 1066
rect -404 678 -346 690
rect -306 1066 -248 1078
rect -306 690 -294 1066
rect -260 690 -248 1066
rect -306 678 -248 690
rect -208 1066 -150 1078
rect -208 690 -196 1066
rect -162 690 -150 1066
rect -208 678 -150 690
rect -110 1066 -52 1078
rect -110 690 -98 1066
rect -64 690 -52 1066
rect -110 678 -52 690
rect -12 1066 46 1078
rect -12 690 0 1066
rect 34 690 46 1066
rect -12 678 46 690
rect 86 1066 144 1078
rect 86 690 98 1066
rect 132 690 144 1066
rect 86 678 144 690
rect 184 1066 242 1078
rect 184 690 196 1066
rect 230 690 242 1066
rect 184 678 242 690
rect 282 1066 340 1078
rect 282 690 294 1066
rect 328 690 340 1066
rect 282 678 340 690
rect 380 1066 438 1078
rect 380 690 392 1066
rect 426 690 438 1066
rect 380 678 438 690
rect 478 1066 536 1078
rect 478 690 490 1066
rect 524 690 536 1066
rect 478 678 536 690
rect 576 1066 634 1078
rect 576 690 588 1066
rect 622 690 634 1066
rect 576 678 634 690
rect 674 1066 732 1078
rect 674 690 686 1066
rect 720 690 732 1066
rect 674 678 732 690
rect 772 1066 830 1078
rect 772 690 784 1066
rect 818 690 830 1066
rect 772 678 830 690
rect 870 1066 928 1078
rect 870 690 882 1066
rect 916 690 928 1066
rect 870 678 928 690
rect 968 1066 1026 1078
rect 968 690 980 1066
rect 1014 690 1026 1066
rect 968 678 1026 690
rect 1066 1066 1124 1078
rect 1066 690 1078 1066
rect 1112 690 1124 1066
rect 1066 678 1124 690
rect 1164 1066 1222 1078
rect 1164 690 1176 1066
rect 1210 690 1222 1066
rect 1164 678 1222 690
rect 1262 1066 1320 1078
rect 1262 690 1274 1066
rect 1308 690 1320 1066
rect 1262 678 1320 690
rect -1188 448 -1130 460
rect -1188 72 -1176 448
rect -1142 72 -1130 448
rect -1188 60 -1130 72
rect -1090 448 -1032 460
rect -1090 72 -1078 448
rect -1044 72 -1032 448
rect -1090 60 -1032 72
rect -992 448 -934 460
rect -992 72 -980 448
rect -946 72 -934 448
rect -992 60 -934 72
rect -894 448 -836 460
rect -894 72 -882 448
rect -848 72 -836 448
rect -894 60 -836 72
rect -796 448 -738 460
rect -796 72 -784 448
rect -750 72 -738 448
rect -796 60 -738 72
rect -698 448 -640 460
rect -698 72 -686 448
rect -652 72 -640 448
rect -698 60 -640 72
rect -600 448 -542 460
rect -600 72 -588 448
rect -554 72 -542 448
rect -600 60 -542 72
rect -502 448 -444 460
rect -502 72 -490 448
rect -456 72 -444 448
rect -502 60 -444 72
rect -404 448 -346 460
rect -404 72 -392 448
rect -358 72 -346 448
rect -404 60 -346 72
rect -306 448 -248 460
rect -306 72 -294 448
rect -260 72 -248 448
rect -306 60 -248 72
rect -208 448 -150 460
rect -208 72 -196 448
rect -162 72 -150 448
rect -208 60 -150 72
rect -110 448 -52 460
rect -110 72 -98 448
rect -64 72 -52 448
rect -110 60 -52 72
rect -12 448 46 460
rect -12 72 0 448
rect 34 72 46 448
rect -12 60 46 72
rect 86 448 144 460
rect 86 72 98 448
rect 132 72 144 448
rect 86 60 144 72
rect 184 448 242 460
rect 184 72 196 448
rect 230 72 242 448
rect 184 60 242 72
rect 282 448 340 460
rect 282 72 294 448
rect 328 72 340 448
rect 282 60 340 72
rect 380 448 438 460
rect 380 72 392 448
rect 426 72 438 448
rect 380 60 438 72
rect 478 448 536 460
rect 478 72 490 448
rect 524 72 536 448
rect 478 60 536 72
rect 576 448 634 460
rect 576 72 588 448
rect 622 72 634 448
rect 576 60 634 72
rect 674 448 732 460
rect 674 72 686 448
rect 720 72 732 448
rect 674 60 732 72
rect 772 448 830 460
rect 772 72 784 448
rect 818 72 830 448
rect 772 60 830 72
rect 870 448 928 460
rect 870 72 882 448
rect 916 72 928 448
rect 870 60 928 72
rect 968 448 1026 460
rect 968 72 980 448
rect 1014 72 1026 448
rect 968 60 1026 72
rect 1066 448 1124 460
rect 1066 72 1078 448
rect 1112 72 1124 448
rect 1066 60 1124 72
rect 1164 448 1222 460
rect 1164 72 1176 448
rect 1210 72 1222 448
rect 1164 60 1222 72
rect 1262 448 1320 460
rect 1262 72 1274 448
rect 1308 72 1320 448
rect 1262 60 1320 72
rect -1188 -378 -1130 -366
rect -1188 -754 -1176 -378
rect -1142 -754 -1130 -378
rect -1188 -766 -1130 -754
rect -1090 -378 -1032 -366
rect -1090 -754 -1078 -378
rect -1044 -754 -1032 -378
rect -1090 -766 -1032 -754
rect -992 -378 -934 -366
rect -992 -754 -980 -378
rect -946 -754 -934 -378
rect -992 -766 -934 -754
rect -894 -378 -836 -366
rect -894 -754 -882 -378
rect -848 -754 -836 -378
rect -894 -766 -836 -754
rect -796 -378 -738 -366
rect -796 -754 -784 -378
rect -750 -754 -738 -378
rect -796 -766 -738 -754
rect -698 -378 -640 -366
rect -698 -754 -686 -378
rect -652 -754 -640 -378
rect -698 -766 -640 -754
rect -600 -378 -542 -366
rect -600 -754 -588 -378
rect -554 -754 -542 -378
rect -600 -766 -542 -754
rect -502 -378 -444 -366
rect -502 -754 -490 -378
rect -456 -754 -444 -378
rect -502 -766 -444 -754
rect -404 -378 -346 -366
rect -404 -754 -392 -378
rect -358 -754 -346 -378
rect -404 -766 -346 -754
rect -306 -378 -248 -366
rect -306 -754 -294 -378
rect -260 -754 -248 -378
rect -306 -766 -248 -754
rect -208 -378 -150 -366
rect -208 -754 -196 -378
rect -162 -754 -150 -378
rect -208 -766 -150 -754
rect -110 -378 -52 -366
rect -110 -754 -98 -378
rect -64 -754 -52 -378
rect -110 -766 -52 -754
rect -12 -378 46 -366
rect -12 -754 0 -378
rect 34 -754 46 -378
rect -12 -766 46 -754
rect 86 -378 144 -366
rect 86 -754 98 -378
rect 132 -754 144 -378
rect 86 -766 144 -754
rect 184 -378 242 -366
rect 184 -754 196 -378
rect 230 -754 242 -378
rect 184 -766 242 -754
rect 282 -378 340 -366
rect 282 -754 294 -378
rect 328 -754 340 -378
rect 282 -766 340 -754
rect 380 -378 438 -366
rect 380 -754 392 -378
rect 426 -754 438 -378
rect 380 -766 438 -754
rect 478 -378 536 -366
rect 478 -754 490 -378
rect 524 -754 536 -378
rect 478 -766 536 -754
rect 576 -378 634 -366
rect 576 -754 588 -378
rect 622 -754 634 -378
rect 576 -766 634 -754
rect 674 -378 732 -366
rect 674 -754 686 -378
rect 720 -754 732 -378
rect 674 -766 732 -754
rect 772 -378 830 -366
rect 772 -754 784 -378
rect 818 -754 830 -378
rect 772 -766 830 -754
rect 870 -378 928 -366
rect 870 -754 882 -378
rect 916 -754 928 -378
rect 870 -766 928 -754
rect 968 -378 1026 -366
rect 968 -754 980 -378
rect 1014 -754 1026 -378
rect 968 -766 1026 -754
rect 1066 -378 1124 -366
rect 1066 -754 1078 -378
rect 1112 -754 1124 -378
rect 1066 -766 1124 -754
rect 1164 -378 1222 -366
rect 1164 -754 1176 -378
rect 1210 -754 1222 -378
rect 1164 -766 1222 -754
rect 1262 -378 1320 -366
rect 1262 -754 1274 -378
rect 1308 -754 1320 -378
rect 1262 -766 1320 -754
rect -1188 -996 -1130 -984
rect -1188 -1372 -1176 -996
rect -1142 -1372 -1130 -996
rect -1188 -1384 -1130 -1372
rect -1090 -996 -1032 -984
rect -1090 -1372 -1078 -996
rect -1044 -1372 -1032 -996
rect -1090 -1384 -1032 -1372
rect -992 -996 -934 -984
rect -992 -1372 -980 -996
rect -946 -1372 -934 -996
rect -992 -1384 -934 -1372
rect -894 -996 -836 -984
rect -894 -1372 -882 -996
rect -848 -1372 -836 -996
rect -894 -1384 -836 -1372
rect -796 -996 -738 -984
rect -796 -1372 -784 -996
rect -750 -1372 -738 -996
rect -796 -1384 -738 -1372
rect -698 -996 -640 -984
rect -698 -1372 -686 -996
rect -652 -1372 -640 -996
rect -698 -1384 -640 -1372
rect -600 -996 -542 -984
rect -600 -1372 -588 -996
rect -554 -1372 -542 -996
rect -600 -1384 -542 -1372
rect -502 -996 -444 -984
rect -502 -1372 -490 -996
rect -456 -1372 -444 -996
rect -502 -1384 -444 -1372
rect -404 -996 -346 -984
rect -404 -1372 -392 -996
rect -358 -1372 -346 -996
rect -404 -1384 -346 -1372
rect -306 -996 -248 -984
rect -306 -1372 -294 -996
rect -260 -1372 -248 -996
rect -306 -1384 -248 -1372
rect -208 -996 -150 -984
rect -208 -1372 -196 -996
rect -162 -1372 -150 -996
rect -208 -1384 -150 -1372
rect -110 -996 -52 -984
rect -110 -1372 -98 -996
rect -64 -1372 -52 -996
rect -110 -1384 -52 -1372
rect -12 -996 46 -984
rect -12 -1372 0 -996
rect 34 -1372 46 -996
rect -12 -1384 46 -1372
rect 86 -996 144 -984
rect 86 -1372 98 -996
rect 132 -1372 144 -996
rect 86 -1384 144 -1372
rect 184 -996 242 -984
rect 184 -1372 196 -996
rect 230 -1372 242 -996
rect 184 -1384 242 -1372
rect 282 -996 340 -984
rect 282 -1372 294 -996
rect 328 -1372 340 -996
rect 282 -1384 340 -1372
rect 380 -996 438 -984
rect 380 -1372 392 -996
rect 426 -1372 438 -996
rect 380 -1384 438 -1372
rect 478 -996 536 -984
rect 478 -1372 490 -996
rect 524 -1372 536 -996
rect 478 -1384 536 -1372
rect 576 -996 634 -984
rect 576 -1372 588 -996
rect 622 -1372 634 -996
rect 576 -1384 634 -1372
rect 674 -996 732 -984
rect 674 -1372 686 -996
rect 720 -1372 732 -996
rect 674 -1384 732 -1372
rect 772 -996 830 -984
rect 772 -1372 784 -996
rect 818 -1372 830 -996
rect 772 -1384 830 -1372
rect 870 -996 928 -984
rect 870 -1372 882 -996
rect 916 -1372 928 -996
rect 870 -1384 928 -1372
rect 968 -996 1026 -984
rect 968 -1372 980 -996
rect 1014 -1372 1026 -996
rect 968 -1384 1026 -1372
rect 1066 -996 1124 -984
rect 1066 -1372 1078 -996
rect 1112 -1372 1124 -996
rect 1066 -1384 1124 -1372
rect 1164 -996 1222 -984
rect 1164 -1372 1176 -996
rect 1210 -1372 1222 -996
rect 1164 -1384 1222 -1372
rect 1262 -996 1320 -984
rect 1262 -1372 1274 -996
rect 1308 -1372 1320 -996
rect 1262 -1384 1320 -1372
rect 2472 746 2530 758
rect 2472 370 2484 746
rect 2518 370 2530 746
rect 2472 358 2530 370
rect 2570 746 2628 758
rect 2570 370 2582 746
rect 2616 370 2628 746
rect 2570 358 2628 370
rect 2668 746 2726 758
rect 2668 370 2680 746
rect 2714 370 2726 746
rect 2668 358 2726 370
rect 2766 746 2824 758
rect 2766 370 2778 746
rect 2812 370 2824 746
rect 2766 358 2824 370
rect 2864 746 2922 758
rect 2864 370 2876 746
rect 2910 370 2922 746
rect 2864 358 2922 370
rect 2962 746 3020 758
rect 2962 370 2974 746
rect 3008 370 3020 746
rect 2962 358 3020 370
rect 3060 746 3118 758
rect 3060 370 3072 746
rect 3106 370 3118 746
rect 3060 358 3118 370
rect 3158 746 3216 758
rect 3158 370 3170 746
rect 3204 370 3216 746
rect 3158 358 3216 370
rect 3256 746 3314 758
rect 3256 370 3268 746
rect 3302 370 3314 746
rect 3256 358 3314 370
rect 3354 746 3412 758
rect 3354 370 3366 746
rect 3400 370 3412 746
rect 3354 358 3412 370
rect 3452 746 3510 758
rect 3452 370 3464 746
rect 3498 370 3510 746
rect 3452 358 3510 370
rect 3550 746 3608 758
rect 3550 370 3562 746
rect 3596 370 3608 746
rect 3550 358 3608 370
rect 3648 746 3706 758
rect 3648 370 3660 746
rect 3694 370 3706 746
rect 3648 358 3706 370
rect 3746 746 3804 758
rect 3746 370 3758 746
rect 3792 370 3804 746
rect 3746 358 3804 370
rect 3844 746 3902 758
rect 3844 370 3856 746
rect 3890 370 3902 746
rect 3844 358 3902 370
rect 3942 746 4000 758
rect 3942 370 3954 746
rect 3988 370 4000 746
rect 3942 358 4000 370
rect 2472 128 2530 140
rect 2472 -248 2484 128
rect 2518 -248 2530 128
rect 2472 -260 2530 -248
rect 2570 128 2628 140
rect 2570 -248 2582 128
rect 2616 -248 2628 128
rect 2570 -260 2628 -248
rect 2668 128 2726 140
rect 2668 -248 2680 128
rect 2714 -248 2726 128
rect 2668 -260 2726 -248
rect 2766 128 2824 140
rect 2766 -248 2778 128
rect 2812 -248 2824 128
rect 2766 -260 2824 -248
rect 2864 128 2922 140
rect 2864 -248 2876 128
rect 2910 -248 2922 128
rect 2864 -260 2922 -248
rect 2962 128 3020 140
rect 2962 -248 2974 128
rect 3008 -248 3020 128
rect 2962 -260 3020 -248
rect 3060 128 3118 140
rect 3060 -248 3072 128
rect 3106 -248 3118 128
rect 3060 -260 3118 -248
rect 3158 128 3216 140
rect 3158 -248 3170 128
rect 3204 -248 3216 128
rect 3158 -260 3216 -248
rect 3256 128 3314 140
rect 3256 -248 3268 128
rect 3302 -248 3314 128
rect 3256 -260 3314 -248
rect 3354 128 3412 140
rect 3354 -248 3366 128
rect 3400 -248 3412 128
rect 3354 -260 3412 -248
rect 3452 128 3510 140
rect 3452 -248 3464 128
rect 3498 -248 3510 128
rect 3452 -260 3510 -248
rect 3550 128 3608 140
rect 3550 -248 3562 128
rect 3596 -248 3608 128
rect 3550 -260 3608 -248
rect 3648 128 3706 140
rect 3648 -248 3660 128
rect 3694 -248 3706 128
rect 3648 -260 3706 -248
rect 3746 128 3804 140
rect 3746 -248 3758 128
rect 3792 -248 3804 128
rect 3746 -260 3804 -248
rect 3844 128 3902 140
rect 3844 -248 3856 128
rect 3890 -248 3902 128
rect 3844 -260 3902 -248
rect 3942 128 4000 140
rect 3942 -248 3954 128
rect 3988 -248 4000 128
rect 3942 -260 4000 -248
rect 1602 -1032 1664 -1020
rect 1602 -1408 1614 -1032
rect 1648 -1408 1664 -1032
rect 1602 -1420 1664 -1408
rect 1694 -1032 1760 -1020
rect 1694 -1408 1710 -1032
rect 1744 -1408 1760 -1032
rect 1694 -1420 1760 -1408
rect 1790 -1032 1856 -1020
rect 1790 -1408 1806 -1032
rect 1840 -1408 1856 -1032
rect 1790 -1420 1856 -1408
rect 1886 -1032 1952 -1020
rect 1886 -1408 1902 -1032
rect 1936 -1408 1952 -1032
rect 1886 -1420 1952 -1408
rect 1982 -1032 2048 -1020
rect 1982 -1408 1998 -1032
rect 2032 -1408 2048 -1032
rect 1982 -1420 2048 -1408
rect 2078 -1032 2144 -1020
rect 2078 -1408 2094 -1032
rect 2128 -1408 2144 -1032
rect 2078 -1420 2144 -1408
rect 2174 -1032 2240 -1020
rect 2174 -1408 2190 -1032
rect 2224 -1408 2240 -1032
rect 2174 -1420 2240 -1408
rect 2270 -1032 2336 -1020
rect 2270 -1408 2286 -1032
rect 2320 -1408 2336 -1032
rect 2270 -1420 2336 -1408
rect 2366 -1032 2432 -1020
rect 2366 -1408 2382 -1032
rect 2416 -1408 2432 -1032
rect 2366 -1420 2432 -1408
rect 2462 -1032 2528 -1020
rect 2462 -1408 2478 -1032
rect 2512 -1408 2528 -1032
rect 2462 -1420 2528 -1408
rect 2558 -1032 2624 -1020
rect 2558 -1408 2574 -1032
rect 2608 -1408 2624 -1032
rect 2558 -1420 2624 -1408
rect 2654 -1032 2720 -1020
rect 2654 -1408 2670 -1032
rect 2704 -1408 2720 -1032
rect 2654 -1420 2720 -1408
rect 2750 -1032 2812 -1020
rect 2750 -1408 2766 -1032
rect 2800 -1408 2812 -1032
rect 2750 -1420 2812 -1408
rect -1208 -1798 -1146 -1786
rect -1208 -2174 -1196 -1798
rect -1162 -2174 -1146 -1798
rect -1208 -2186 -1146 -2174
rect -1116 -1798 -1050 -1786
rect -1116 -2174 -1100 -1798
rect -1066 -2174 -1050 -1798
rect -1116 -2186 -1050 -2174
rect -1020 -1798 -954 -1786
rect -1020 -2174 -1004 -1798
rect -970 -2174 -954 -1798
rect -1020 -2186 -954 -2174
rect -924 -1798 -858 -1786
rect -924 -2174 -908 -1798
rect -874 -2174 -858 -1798
rect -924 -2186 -858 -2174
rect -828 -1798 -762 -1786
rect -828 -2174 -812 -1798
rect -778 -2174 -762 -1798
rect -828 -2186 -762 -2174
rect -732 -1798 -666 -1786
rect -732 -2174 -716 -1798
rect -682 -2174 -666 -1798
rect -732 -2186 -666 -2174
rect -636 -1798 -570 -1786
rect -636 -2174 -620 -1798
rect -586 -2174 -570 -1798
rect -636 -2186 -570 -2174
rect -540 -1798 -474 -1786
rect -540 -2174 -524 -1798
rect -490 -2174 -474 -1798
rect -540 -2186 -474 -2174
rect -444 -1798 -378 -1786
rect -444 -2174 -428 -1798
rect -394 -2174 -378 -1798
rect -444 -2186 -378 -2174
rect -348 -1798 -282 -1786
rect -348 -2174 -332 -1798
rect -298 -2174 -282 -1798
rect -348 -2186 -282 -2174
rect -252 -1798 -186 -1786
rect -252 -2174 -236 -1798
rect -202 -2174 -186 -1798
rect -252 -2186 -186 -2174
rect -156 -1798 -90 -1786
rect -156 -2174 -140 -1798
rect -106 -2174 -90 -1798
rect -156 -2186 -90 -2174
rect -60 -1798 6 -1786
rect -60 -2174 -44 -1798
rect -10 -2174 6 -1798
rect -60 -2186 6 -2174
rect 36 -1798 102 -1786
rect 36 -2174 52 -1798
rect 86 -2174 102 -1798
rect 36 -2186 102 -2174
rect 132 -1798 198 -1786
rect 132 -2174 148 -1798
rect 182 -2174 198 -1798
rect 132 -2186 198 -2174
rect 228 -1798 294 -1786
rect 228 -2174 244 -1798
rect 278 -2174 294 -1798
rect 228 -2186 294 -2174
rect 324 -1798 390 -1786
rect 324 -2174 340 -1798
rect 374 -2174 390 -1798
rect 324 -2186 390 -2174
rect 420 -1798 486 -1786
rect 420 -2174 436 -1798
rect 470 -2174 486 -1798
rect 420 -2186 486 -2174
rect 516 -1798 582 -1786
rect 516 -2174 532 -1798
rect 566 -2174 582 -1798
rect 516 -2186 582 -2174
rect 612 -1798 678 -1786
rect 612 -2174 628 -1798
rect 662 -2174 678 -1798
rect 612 -2186 678 -2174
rect 708 -1798 774 -1786
rect 708 -2174 724 -1798
rect 758 -2174 774 -1798
rect 708 -2186 774 -2174
rect 804 -1798 870 -1786
rect 804 -2174 820 -1798
rect 854 -2174 870 -1798
rect 804 -2186 870 -2174
rect 900 -1798 966 -1786
rect 900 -2174 916 -1798
rect 950 -2174 966 -1798
rect 900 -2186 966 -2174
rect 996 -1798 1062 -1786
rect 996 -2174 1012 -1798
rect 1046 -2174 1062 -1798
rect 996 -2186 1062 -2174
rect 1092 -1798 1158 -1786
rect 1092 -2174 1108 -1798
rect 1142 -2174 1158 -1798
rect 1092 -2186 1158 -2174
rect 1188 -1798 1250 -1786
rect 1188 -2174 1204 -1798
rect 1238 -2174 1250 -1798
rect 1188 -2186 1250 -2174
rect -1208 -2416 -1146 -2404
rect -1208 -2792 -1196 -2416
rect -1162 -2792 -1146 -2416
rect -1208 -2804 -1146 -2792
rect -1116 -2416 -1050 -2404
rect -1116 -2792 -1100 -2416
rect -1066 -2792 -1050 -2416
rect -1116 -2804 -1050 -2792
rect -1020 -2416 -954 -2404
rect -1020 -2792 -1004 -2416
rect -970 -2792 -954 -2416
rect -1020 -2804 -954 -2792
rect -924 -2416 -858 -2404
rect -924 -2792 -908 -2416
rect -874 -2792 -858 -2416
rect -924 -2804 -858 -2792
rect -828 -2416 -762 -2404
rect -828 -2792 -812 -2416
rect -778 -2792 -762 -2416
rect -828 -2804 -762 -2792
rect -732 -2416 -666 -2404
rect -732 -2792 -716 -2416
rect -682 -2792 -666 -2416
rect -732 -2804 -666 -2792
rect -636 -2416 -570 -2404
rect -636 -2792 -620 -2416
rect -586 -2792 -570 -2416
rect -636 -2804 -570 -2792
rect -540 -2416 -474 -2404
rect -540 -2792 -524 -2416
rect -490 -2792 -474 -2416
rect -540 -2804 -474 -2792
rect -444 -2416 -378 -2404
rect -444 -2792 -428 -2416
rect -394 -2792 -378 -2416
rect -444 -2804 -378 -2792
rect -348 -2416 -282 -2404
rect -348 -2792 -332 -2416
rect -298 -2792 -282 -2416
rect -348 -2804 -282 -2792
rect -252 -2416 -186 -2404
rect -252 -2792 -236 -2416
rect -202 -2792 -186 -2416
rect -252 -2804 -186 -2792
rect -156 -2416 -90 -2404
rect -156 -2792 -140 -2416
rect -106 -2792 -90 -2416
rect -156 -2804 -90 -2792
rect -60 -2416 6 -2404
rect -60 -2792 -44 -2416
rect -10 -2792 6 -2416
rect -60 -2804 6 -2792
rect 36 -2416 102 -2404
rect 36 -2792 52 -2416
rect 86 -2792 102 -2416
rect 36 -2804 102 -2792
rect 132 -2416 198 -2404
rect 132 -2792 148 -2416
rect 182 -2792 198 -2416
rect 132 -2804 198 -2792
rect 228 -2416 294 -2404
rect 228 -2792 244 -2416
rect 278 -2792 294 -2416
rect 228 -2804 294 -2792
rect 324 -2416 390 -2404
rect 324 -2792 340 -2416
rect 374 -2792 390 -2416
rect 324 -2804 390 -2792
rect 420 -2416 486 -2404
rect 420 -2792 436 -2416
rect 470 -2792 486 -2416
rect 420 -2804 486 -2792
rect 516 -2416 582 -2404
rect 516 -2792 532 -2416
rect 566 -2792 582 -2416
rect 516 -2804 582 -2792
rect 612 -2416 678 -2404
rect 612 -2792 628 -2416
rect 662 -2792 678 -2416
rect 612 -2804 678 -2792
rect 708 -2416 774 -2404
rect 708 -2792 724 -2416
rect 758 -2792 774 -2416
rect 708 -2804 774 -2792
rect 804 -2416 870 -2404
rect 804 -2792 820 -2416
rect 854 -2792 870 -2416
rect 804 -2804 870 -2792
rect 900 -2416 966 -2404
rect 900 -2792 916 -2416
rect 950 -2792 966 -2416
rect 900 -2804 966 -2792
rect 996 -2416 1062 -2404
rect 996 -2792 1012 -2416
rect 1046 -2792 1062 -2416
rect 996 -2804 1062 -2792
rect 1092 -2416 1158 -2404
rect 1092 -2792 1108 -2416
rect 1142 -2792 1158 -2416
rect 1092 -2804 1158 -2792
rect 1188 -2416 1250 -2404
rect 1188 -2792 1204 -2416
rect 1238 -2792 1250 -2416
rect 1188 -2804 1250 -2792
rect -1208 -3034 -1146 -3022
rect -1208 -3410 -1196 -3034
rect -1162 -3410 -1146 -3034
rect -1208 -3422 -1146 -3410
rect -1116 -3034 -1050 -3022
rect -1116 -3410 -1100 -3034
rect -1066 -3410 -1050 -3034
rect -1116 -3422 -1050 -3410
rect -1020 -3034 -954 -3022
rect -1020 -3410 -1004 -3034
rect -970 -3410 -954 -3034
rect -1020 -3422 -954 -3410
rect -924 -3034 -858 -3022
rect -924 -3410 -908 -3034
rect -874 -3410 -858 -3034
rect -924 -3422 -858 -3410
rect -828 -3034 -762 -3022
rect -828 -3410 -812 -3034
rect -778 -3410 -762 -3034
rect -828 -3422 -762 -3410
rect -732 -3034 -666 -3022
rect -732 -3410 -716 -3034
rect -682 -3410 -666 -3034
rect -732 -3422 -666 -3410
rect -636 -3034 -570 -3022
rect -636 -3410 -620 -3034
rect -586 -3410 -570 -3034
rect -636 -3422 -570 -3410
rect -540 -3034 -474 -3022
rect -540 -3410 -524 -3034
rect -490 -3410 -474 -3034
rect -540 -3422 -474 -3410
rect -444 -3034 -378 -3022
rect -444 -3410 -428 -3034
rect -394 -3410 -378 -3034
rect -444 -3422 -378 -3410
rect -348 -3034 -282 -3022
rect -348 -3410 -332 -3034
rect -298 -3410 -282 -3034
rect -348 -3422 -282 -3410
rect -252 -3034 -186 -3022
rect -252 -3410 -236 -3034
rect -202 -3410 -186 -3034
rect -252 -3422 -186 -3410
rect -156 -3034 -90 -3022
rect -156 -3410 -140 -3034
rect -106 -3410 -90 -3034
rect -156 -3422 -90 -3410
rect -60 -3034 6 -3022
rect -60 -3410 -44 -3034
rect -10 -3410 6 -3034
rect -60 -3422 6 -3410
rect 36 -3034 102 -3022
rect 36 -3410 52 -3034
rect 86 -3410 102 -3034
rect 36 -3422 102 -3410
rect 132 -3034 198 -3022
rect 132 -3410 148 -3034
rect 182 -3410 198 -3034
rect 132 -3422 198 -3410
rect 228 -3034 294 -3022
rect 228 -3410 244 -3034
rect 278 -3410 294 -3034
rect 228 -3422 294 -3410
rect 324 -3034 390 -3022
rect 324 -3410 340 -3034
rect 374 -3410 390 -3034
rect 324 -3422 390 -3410
rect 420 -3034 486 -3022
rect 420 -3410 436 -3034
rect 470 -3410 486 -3034
rect 420 -3422 486 -3410
rect 516 -3034 582 -3022
rect 516 -3410 532 -3034
rect 566 -3410 582 -3034
rect 516 -3422 582 -3410
rect 612 -3034 678 -3022
rect 612 -3410 628 -3034
rect 662 -3410 678 -3034
rect 612 -3422 678 -3410
rect 708 -3034 774 -3022
rect 708 -3410 724 -3034
rect 758 -3410 774 -3034
rect 708 -3422 774 -3410
rect 804 -3034 870 -3022
rect 804 -3410 820 -3034
rect 854 -3410 870 -3034
rect 804 -3422 870 -3410
rect 900 -3034 966 -3022
rect 900 -3410 916 -3034
rect 950 -3410 966 -3034
rect 900 -3422 966 -3410
rect 996 -3034 1062 -3022
rect 996 -3410 1012 -3034
rect 1046 -3410 1062 -3034
rect 996 -3422 1062 -3410
rect 1092 -3034 1158 -3022
rect 1092 -3410 1108 -3034
rect 1142 -3410 1158 -3034
rect 1092 -3422 1158 -3410
rect 1188 -3034 1250 -3022
rect 1188 -3410 1204 -3034
rect 1238 -3410 1250 -3034
rect 1188 -3422 1250 -3410
rect -1208 -3652 -1146 -3640
rect -1208 -4028 -1196 -3652
rect -1162 -4028 -1146 -3652
rect -1208 -4040 -1146 -4028
rect -1116 -3652 -1050 -3640
rect -1116 -4028 -1100 -3652
rect -1066 -4028 -1050 -3652
rect -1116 -4040 -1050 -4028
rect -1020 -3652 -954 -3640
rect -1020 -4028 -1004 -3652
rect -970 -4028 -954 -3652
rect -1020 -4040 -954 -4028
rect -924 -3652 -858 -3640
rect -924 -4028 -908 -3652
rect -874 -4028 -858 -3652
rect -924 -4040 -858 -4028
rect -828 -3652 -762 -3640
rect -828 -4028 -812 -3652
rect -778 -4028 -762 -3652
rect -828 -4040 -762 -4028
rect -732 -3652 -666 -3640
rect -732 -4028 -716 -3652
rect -682 -4028 -666 -3652
rect -732 -4040 -666 -4028
rect -636 -3652 -570 -3640
rect -636 -4028 -620 -3652
rect -586 -4028 -570 -3652
rect -636 -4040 -570 -4028
rect -540 -3652 -474 -3640
rect -540 -4028 -524 -3652
rect -490 -4028 -474 -3652
rect -540 -4040 -474 -4028
rect -444 -3652 -378 -3640
rect -444 -4028 -428 -3652
rect -394 -4028 -378 -3652
rect -444 -4040 -378 -4028
rect -348 -3652 -282 -3640
rect -348 -4028 -332 -3652
rect -298 -4028 -282 -3652
rect -348 -4040 -282 -4028
rect -252 -3652 -186 -3640
rect -252 -4028 -236 -3652
rect -202 -4028 -186 -3652
rect -252 -4040 -186 -4028
rect -156 -3652 -90 -3640
rect -156 -4028 -140 -3652
rect -106 -4028 -90 -3652
rect -156 -4040 -90 -4028
rect -60 -3652 6 -3640
rect -60 -4028 -44 -3652
rect -10 -4028 6 -3652
rect -60 -4040 6 -4028
rect 36 -3652 102 -3640
rect 36 -4028 52 -3652
rect 86 -4028 102 -3652
rect 36 -4040 102 -4028
rect 132 -3652 198 -3640
rect 132 -4028 148 -3652
rect 182 -4028 198 -3652
rect 132 -4040 198 -4028
rect 228 -3652 294 -3640
rect 228 -4028 244 -3652
rect 278 -4028 294 -3652
rect 228 -4040 294 -4028
rect 324 -3652 390 -3640
rect 324 -4028 340 -3652
rect 374 -4028 390 -3652
rect 324 -4040 390 -4028
rect 420 -3652 486 -3640
rect 420 -4028 436 -3652
rect 470 -4028 486 -3652
rect 420 -4040 486 -4028
rect 516 -3652 582 -3640
rect 516 -4028 532 -3652
rect 566 -4028 582 -3652
rect 516 -4040 582 -4028
rect 612 -3652 678 -3640
rect 612 -4028 628 -3652
rect 662 -4028 678 -3652
rect 612 -4040 678 -4028
rect 708 -3652 774 -3640
rect 708 -4028 724 -3652
rect 758 -4028 774 -3652
rect 708 -4040 774 -4028
rect 804 -3652 870 -3640
rect 804 -4028 820 -3652
rect 854 -4028 870 -3652
rect 804 -4040 870 -4028
rect 900 -3652 966 -3640
rect 900 -4028 916 -3652
rect 950 -4028 966 -3652
rect 900 -4040 966 -4028
rect 996 -3652 1062 -3640
rect 996 -4028 1012 -3652
rect 1046 -4028 1062 -3652
rect 996 -4040 1062 -4028
rect 1092 -3652 1158 -3640
rect 1092 -4028 1108 -3652
rect 1142 -4028 1158 -3652
rect 1092 -4040 1158 -4028
rect 1188 -3652 1250 -3640
rect 1188 -4028 1204 -3652
rect 1238 -4028 1250 -3652
rect 1188 -4040 1250 -4028
rect 1602 -1852 1660 -1840
rect 1602 -2228 1614 -1852
rect 1648 -2228 1660 -1852
rect 1602 -2240 1660 -2228
rect 1860 -1852 1918 -1840
rect 1860 -2228 1872 -1852
rect 1906 -2228 1918 -1852
rect 1860 -2240 1918 -2228
rect 2118 -1852 2176 -1840
rect 2118 -2228 2130 -1852
rect 2164 -2228 2176 -1852
rect 2118 -2240 2176 -2228
rect 2376 -1852 2434 -1840
rect 2376 -2228 2388 -1852
rect 2422 -2228 2434 -1852
rect 2376 -2240 2434 -2228
rect 2634 -1852 2692 -1840
rect 2634 -2228 2646 -1852
rect 2680 -2228 2692 -1852
rect 2634 -2240 2692 -2228
rect 2892 -1852 2950 -1840
rect 2892 -2228 2904 -1852
rect 2938 -2228 2950 -1852
rect 2892 -2240 2950 -2228
rect 3150 -1852 3208 -1840
rect 3150 -2228 3162 -1852
rect 3196 -2228 3208 -1852
rect 3150 -2240 3208 -2228
rect -1188 -6004 -1130 -5992
rect -1188 -6380 -1176 -6004
rect -1142 -6380 -1130 -6004
rect -1188 -6392 -1130 -6380
rect -1090 -6004 -1032 -5992
rect -1090 -6380 -1078 -6004
rect -1044 -6380 -1032 -6004
rect -1090 -6392 -1032 -6380
rect -992 -6004 -934 -5992
rect -992 -6380 -980 -6004
rect -946 -6380 -934 -6004
rect -992 -6392 -934 -6380
rect -894 -6004 -836 -5992
rect -894 -6380 -882 -6004
rect -848 -6380 -836 -6004
rect -894 -6392 -836 -6380
rect -796 -6004 -738 -5992
rect -796 -6380 -784 -6004
rect -750 -6380 -738 -6004
rect -796 -6392 -738 -6380
rect -698 -6004 -640 -5992
rect -698 -6380 -686 -6004
rect -652 -6380 -640 -6004
rect -698 -6392 -640 -6380
rect -600 -6004 -542 -5992
rect -600 -6380 -588 -6004
rect -554 -6380 -542 -6004
rect -600 -6392 -542 -6380
rect -502 -6004 -444 -5992
rect -502 -6380 -490 -6004
rect -456 -6380 -444 -6004
rect -502 -6392 -444 -6380
rect -404 -6004 -346 -5992
rect -404 -6380 -392 -6004
rect -358 -6380 -346 -6004
rect -404 -6392 -346 -6380
rect -306 -6004 -248 -5992
rect -306 -6380 -294 -6004
rect -260 -6380 -248 -6004
rect -306 -6392 -248 -6380
rect -208 -6004 -150 -5992
rect -208 -6380 -196 -6004
rect -162 -6380 -150 -6004
rect -208 -6392 -150 -6380
rect -110 -6004 -52 -5992
rect -110 -6380 -98 -6004
rect -64 -6380 -52 -6004
rect -110 -6392 -52 -6380
rect -12 -6004 46 -5992
rect -12 -6380 0 -6004
rect 34 -6380 46 -6004
rect -12 -6392 46 -6380
rect 86 -6004 144 -5992
rect 86 -6380 98 -6004
rect 132 -6380 144 -6004
rect 86 -6392 144 -6380
rect 184 -6004 242 -5992
rect 184 -6380 196 -6004
rect 230 -6380 242 -6004
rect 184 -6392 242 -6380
rect 282 -6004 340 -5992
rect 282 -6380 294 -6004
rect 328 -6380 340 -6004
rect 282 -6392 340 -6380
rect 380 -6004 438 -5992
rect 380 -6380 392 -6004
rect 426 -6380 438 -6004
rect 380 -6392 438 -6380
rect 478 -6004 536 -5992
rect 478 -6380 490 -6004
rect 524 -6380 536 -6004
rect 478 -6392 536 -6380
rect 576 -6004 634 -5992
rect 576 -6380 588 -6004
rect 622 -6380 634 -6004
rect 576 -6392 634 -6380
rect 674 -6004 732 -5992
rect 674 -6380 686 -6004
rect 720 -6380 732 -6004
rect 674 -6392 732 -6380
rect 772 -6004 830 -5992
rect 772 -6380 784 -6004
rect 818 -6380 830 -6004
rect 772 -6392 830 -6380
rect 870 -6004 928 -5992
rect 870 -6380 882 -6004
rect 916 -6380 928 -6004
rect 870 -6392 928 -6380
rect 968 -6004 1026 -5992
rect 968 -6380 980 -6004
rect 1014 -6380 1026 -6004
rect 968 -6392 1026 -6380
rect 1066 -6004 1124 -5992
rect 1066 -6380 1078 -6004
rect 1112 -6380 1124 -6004
rect 1066 -6392 1124 -6380
rect 1164 -6004 1222 -5992
rect 1164 -6380 1176 -6004
rect 1210 -6380 1222 -6004
rect 1164 -6392 1222 -6380
rect 1262 -6004 1320 -5992
rect 1262 -6380 1274 -6004
rect 1308 -6380 1320 -6004
rect 1262 -6392 1320 -6380
rect -1188 -6622 -1130 -6610
rect -1188 -6998 -1176 -6622
rect -1142 -6998 -1130 -6622
rect -1188 -7010 -1130 -6998
rect -1090 -6622 -1032 -6610
rect -1090 -6998 -1078 -6622
rect -1044 -6998 -1032 -6622
rect -1090 -7010 -1032 -6998
rect -992 -6622 -934 -6610
rect -992 -6998 -980 -6622
rect -946 -6998 -934 -6622
rect -992 -7010 -934 -6998
rect -894 -6622 -836 -6610
rect -894 -6998 -882 -6622
rect -848 -6998 -836 -6622
rect -894 -7010 -836 -6998
rect -796 -6622 -738 -6610
rect -796 -6998 -784 -6622
rect -750 -6998 -738 -6622
rect -796 -7010 -738 -6998
rect -698 -6622 -640 -6610
rect -698 -6998 -686 -6622
rect -652 -6998 -640 -6622
rect -698 -7010 -640 -6998
rect -600 -6622 -542 -6610
rect -600 -6998 -588 -6622
rect -554 -6998 -542 -6622
rect -600 -7010 -542 -6998
rect -502 -6622 -444 -6610
rect -502 -6998 -490 -6622
rect -456 -6998 -444 -6622
rect -502 -7010 -444 -6998
rect -404 -6622 -346 -6610
rect -404 -6998 -392 -6622
rect -358 -6998 -346 -6622
rect -404 -7010 -346 -6998
rect -306 -6622 -248 -6610
rect -306 -6998 -294 -6622
rect -260 -6998 -248 -6622
rect -306 -7010 -248 -6998
rect -208 -6622 -150 -6610
rect -208 -6998 -196 -6622
rect -162 -6998 -150 -6622
rect -208 -7010 -150 -6998
rect -110 -6622 -52 -6610
rect -110 -6998 -98 -6622
rect -64 -6998 -52 -6622
rect -110 -7010 -52 -6998
rect -12 -6622 46 -6610
rect -12 -6998 0 -6622
rect 34 -6998 46 -6622
rect -12 -7010 46 -6998
rect 86 -6622 144 -6610
rect 86 -6998 98 -6622
rect 132 -6998 144 -6622
rect 86 -7010 144 -6998
rect 184 -6622 242 -6610
rect 184 -6998 196 -6622
rect 230 -6998 242 -6622
rect 184 -7010 242 -6998
rect 282 -6622 340 -6610
rect 282 -6998 294 -6622
rect 328 -6998 340 -6622
rect 282 -7010 340 -6998
rect 380 -6622 438 -6610
rect 380 -6998 392 -6622
rect 426 -6998 438 -6622
rect 380 -7010 438 -6998
rect 478 -6622 536 -6610
rect 478 -6998 490 -6622
rect 524 -6998 536 -6622
rect 478 -7010 536 -6998
rect 576 -6622 634 -6610
rect 576 -6998 588 -6622
rect 622 -6998 634 -6622
rect 576 -7010 634 -6998
rect 674 -6622 732 -6610
rect 674 -6998 686 -6622
rect 720 -6998 732 -6622
rect 674 -7010 732 -6998
rect 772 -6622 830 -6610
rect 772 -6998 784 -6622
rect 818 -6998 830 -6622
rect 772 -7010 830 -6998
rect 870 -6622 928 -6610
rect 870 -6998 882 -6622
rect 916 -6998 928 -6622
rect 870 -7010 928 -6998
rect 968 -6622 1026 -6610
rect 968 -6998 980 -6622
rect 1014 -6998 1026 -6622
rect 968 -7010 1026 -6998
rect 1066 -6622 1124 -6610
rect 1066 -6998 1078 -6622
rect 1112 -6998 1124 -6622
rect 1066 -7010 1124 -6998
rect 1164 -6622 1222 -6610
rect 1164 -6998 1176 -6622
rect 1210 -6998 1222 -6622
rect 1164 -7010 1222 -6998
rect 1262 -6622 1320 -6610
rect 1262 -6998 1274 -6622
rect 1308 -6998 1320 -6622
rect 1262 -7010 1320 -6998
rect -1188 -7448 -1130 -7436
rect -1188 -7824 -1176 -7448
rect -1142 -7824 -1130 -7448
rect -1188 -7836 -1130 -7824
rect -1090 -7448 -1032 -7436
rect -1090 -7824 -1078 -7448
rect -1044 -7824 -1032 -7448
rect -1090 -7836 -1032 -7824
rect -992 -7448 -934 -7436
rect -992 -7824 -980 -7448
rect -946 -7824 -934 -7448
rect -992 -7836 -934 -7824
rect -894 -7448 -836 -7436
rect -894 -7824 -882 -7448
rect -848 -7824 -836 -7448
rect -894 -7836 -836 -7824
rect -796 -7448 -738 -7436
rect -796 -7824 -784 -7448
rect -750 -7824 -738 -7448
rect -796 -7836 -738 -7824
rect -698 -7448 -640 -7436
rect -698 -7824 -686 -7448
rect -652 -7824 -640 -7448
rect -698 -7836 -640 -7824
rect -600 -7448 -542 -7436
rect -600 -7824 -588 -7448
rect -554 -7824 -542 -7448
rect -600 -7836 -542 -7824
rect -502 -7448 -444 -7436
rect -502 -7824 -490 -7448
rect -456 -7824 -444 -7448
rect -502 -7836 -444 -7824
rect -404 -7448 -346 -7436
rect -404 -7824 -392 -7448
rect -358 -7824 -346 -7448
rect -404 -7836 -346 -7824
rect -306 -7448 -248 -7436
rect -306 -7824 -294 -7448
rect -260 -7824 -248 -7448
rect -306 -7836 -248 -7824
rect -208 -7448 -150 -7436
rect -208 -7824 -196 -7448
rect -162 -7824 -150 -7448
rect -208 -7836 -150 -7824
rect -110 -7448 -52 -7436
rect -110 -7824 -98 -7448
rect -64 -7824 -52 -7448
rect -110 -7836 -52 -7824
rect -12 -7448 46 -7436
rect -12 -7824 0 -7448
rect 34 -7824 46 -7448
rect -12 -7836 46 -7824
rect 86 -7448 144 -7436
rect 86 -7824 98 -7448
rect 132 -7824 144 -7448
rect 86 -7836 144 -7824
rect 184 -7448 242 -7436
rect 184 -7824 196 -7448
rect 230 -7824 242 -7448
rect 184 -7836 242 -7824
rect 282 -7448 340 -7436
rect 282 -7824 294 -7448
rect 328 -7824 340 -7448
rect 282 -7836 340 -7824
rect 380 -7448 438 -7436
rect 380 -7824 392 -7448
rect 426 -7824 438 -7448
rect 380 -7836 438 -7824
rect 478 -7448 536 -7436
rect 478 -7824 490 -7448
rect 524 -7824 536 -7448
rect 478 -7836 536 -7824
rect 576 -7448 634 -7436
rect 576 -7824 588 -7448
rect 622 -7824 634 -7448
rect 576 -7836 634 -7824
rect 674 -7448 732 -7436
rect 674 -7824 686 -7448
rect 720 -7824 732 -7448
rect 674 -7836 732 -7824
rect 772 -7448 830 -7436
rect 772 -7824 784 -7448
rect 818 -7824 830 -7448
rect 772 -7836 830 -7824
rect 870 -7448 928 -7436
rect 870 -7824 882 -7448
rect 916 -7824 928 -7448
rect 870 -7836 928 -7824
rect 968 -7448 1026 -7436
rect 968 -7824 980 -7448
rect 1014 -7824 1026 -7448
rect 968 -7836 1026 -7824
rect 1066 -7448 1124 -7436
rect 1066 -7824 1078 -7448
rect 1112 -7824 1124 -7448
rect 1066 -7836 1124 -7824
rect 1164 -7448 1222 -7436
rect 1164 -7824 1176 -7448
rect 1210 -7824 1222 -7448
rect 1164 -7836 1222 -7824
rect 1262 -7448 1320 -7436
rect 1262 -7824 1274 -7448
rect 1308 -7824 1320 -7448
rect 1262 -7836 1320 -7824
rect -1188 -8066 -1130 -8054
rect -1188 -8442 -1176 -8066
rect -1142 -8442 -1130 -8066
rect -1188 -8454 -1130 -8442
rect -1090 -8066 -1032 -8054
rect -1090 -8442 -1078 -8066
rect -1044 -8442 -1032 -8066
rect -1090 -8454 -1032 -8442
rect -992 -8066 -934 -8054
rect -992 -8442 -980 -8066
rect -946 -8442 -934 -8066
rect -992 -8454 -934 -8442
rect -894 -8066 -836 -8054
rect -894 -8442 -882 -8066
rect -848 -8442 -836 -8066
rect -894 -8454 -836 -8442
rect -796 -8066 -738 -8054
rect -796 -8442 -784 -8066
rect -750 -8442 -738 -8066
rect -796 -8454 -738 -8442
rect -698 -8066 -640 -8054
rect -698 -8442 -686 -8066
rect -652 -8442 -640 -8066
rect -698 -8454 -640 -8442
rect -600 -8066 -542 -8054
rect -600 -8442 -588 -8066
rect -554 -8442 -542 -8066
rect -600 -8454 -542 -8442
rect -502 -8066 -444 -8054
rect -502 -8442 -490 -8066
rect -456 -8442 -444 -8066
rect -502 -8454 -444 -8442
rect -404 -8066 -346 -8054
rect -404 -8442 -392 -8066
rect -358 -8442 -346 -8066
rect -404 -8454 -346 -8442
rect -306 -8066 -248 -8054
rect -306 -8442 -294 -8066
rect -260 -8442 -248 -8066
rect -306 -8454 -248 -8442
rect -208 -8066 -150 -8054
rect -208 -8442 -196 -8066
rect -162 -8442 -150 -8066
rect -208 -8454 -150 -8442
rect -110 -8066 -52 -8054
rect -110 -8442 -98 -8066
rect -64 -8442 -52 -8066
rect -110 -8454 -52 -8442
rect -12 -8066 46 -8054
rect -12 -8442 0 -8066
rect 34 -8442 46 -8066
rect -12 -8454 46 -8442
rect 86 -8066 144 -8054
rect 86 -8442 98 -8066
rect 132 -8442 144 -8066
rect 86 -8454 144 -8442
rect 184 -8066 242 -8054
rect 184 -8442 196 -8066
rect 230 -8442 242 -8066
rect 184 -8454 242 -8442
rect 282 -8066 340 -8054
rect 282 -8442 294 -8066
rect 328 -8442 340 -8066
rect 282 -8454 340 -8442
rect 380 -8066 438 -8054
rect 380 -8442 392 -8066
rect 426 -8442 438 -8066
rect 380 -8454 438 -8442
rect 478 -8066 536 -8054
rect 478 -8442 490 -8066
rect 524 -8442 536 -8066
rect 478 -8454 536 -8442
rect 576 -8066 634 -8054
rect 576 -8442 588 -8066
rect 622 -8442 634 -8066
rect 576 -8454 634 -8442
rect 674 -8066 732 -8054
rect 674 -8442 686 -8066
rect 720 -8442 732 -8066
rect 674 -8454 732 -8442
rect 772 -8066 830 -8054
rect 772 -8442 784 -8066
rect 818 -8442 830 -8066
rect 772 -8454 830 -8442
rect 870 -8066 928 -8054
rect 870 -8442 882 -8066
rect 916 -8442 928 -8066
rect 870 -8454 928 -8442
rect 968 -8066 1026 -8054
rect 968 -8442 980 -8066
rect 1014 -8442 1026 -8066
rect 968 -8454 1026 -8442
rect 1066 -8066 1124 -8054
rect 1066 -8442 1078 -8066
rect 1112 -8442 1124 -8066
rect 1066 -8454 1124 -8442
rect 1164 -8066 1222 -8054
rect 1164 -8442 1176 -8066
rect 1210 -8442 1222 -8066
rect 1164 -8454 1222 -8442
rect 1262 -8066 1320 -8054
rect 1262 -8442 1274 -8066
rect 1308 -8442 1320 -8066
rect 1262 -8454 1320 -8442
rect 2472 -6324 2530 -6312
rect 2472 -6700 2484 -6324
rect 2518 -6700 2530 -6324
rect 2472 -6712 2530 -6700
rect 2570 -6324 2628 -6312
rect 2570 -6700 2582 -6324
rect 2616 -6700 2628 -6324
rect 2570 -6712 2628 -6700
rect 2668 -6324 2726 -6312
rect 2668 -6700 2680 -6324
rect 2714 -6700 2726 -6324
rect 2668 -6712 2726 -6700
rect 2766 -6324 2824 -6312
rect 2766 -6700 2778 -6324
rect 2812 -6700 2824 -6324
rect 2766 -6712 2824 -6700
rect 2864 -6324 2922 -6312
rect 2864 -6700 2876 -6324
rect 2910 -6700 2922 -6324
rect 2864 -6712 2922 -6700
rect 2962 -6324 3020 -6312
rect 2962 -6700 2974 -6324
rect 3008 -6700 3020 -6324
rect 2962 -6712 3020 -6700
rect 3060 -6324 3118 -6312
rect 3060 -6700 3072 -6324
rect 3106 -6700 3118 -6324
rect 3060 -6712 3118 -6700
rect 3158 -6324 3216 -6312
rect 3158 -6700 3170 -6324
rect 3204 -6700 3216 -6324
rect 3158 -6712 3216 -6700
rect 3256 -6324 3314 -6312
rect 3256 -6700 3268 -6324
rect 3302 -6700 3314 -6324
rect 3256 -6712 3314 -6700
rect 3354 -6324 3412 -6312
rect 3354 -6700 3366 -6324
rect 3400 -6700 3412 -6324
rect 3354 -6712 3412 -6700
rect 3452 -6324 3510 -6312
rect 3452 -6700 3464 -6324
rect 3498 -6700 3510 -6324
rect 3452 -6712 3510 -6700
rect 3550 -6324 3608 -6312
rect 3550 -6700 3562 -6324
rect 3596 -6700 3608 -6324
rect 3550 -6712 3608 -6700
rect 3648 -6324 3706 -6312
rect 3648 -6700 3660 -6324
rect 3694 -6700 3706 -6324
rect 3648 -6712 3706 -6700
rect 3746 -6324 3804 -6312
rect 3746 -6700 3758 -6324
rect 3792 -6700 3804 -6324
rect 3746 -6712 3804 -6700
rect 3844 -6324 3902 -6312
rect 3844 -6700 3856 -6324
rect 3890 -6700 3902 -6324
rect 3844 -6712 3902 -6700
rect 3942 -6324 4000 -6312
rect 3942 -6700 3954 -6324
rect 3988 -6700 4000 -6324
rect 3942 -6712 4000 -6700
rect 2472 -6942 2530 -6930
rect 2472 -7318 2484 -6942
rect 2518 -7318 2530 -6942
rect 2472 -7330 2530 -7318
rect 2570 -6942 2628 -6930
rect 2570 -7318 2582 -6942
rect 2616 -7318 2628 -6942
rect 2570 -7330 2628 -7318
rect 2668 -6942 2726 -6930
rect 2668 -7318 2680 -6942
rect 2714 -7318 2726 -6942
rect 2668 -7330 2726 -7318
rect 2766 -6942 2824 -6930
rect 2766 -7318 2778 -6942
rect 2812 -7318 2824 -6942
rect 2766 -7330 2824 -7318
rect 2864 -6942 2922 -6930
rect 2864 -7318 2876 -6942
rect 2910 -7318 2922 -6942
rect 2864 -7330 2922 -7318
rect 2962 -6942 3020 -6930
rect 2962 -7318 2974 -6942
rect 3008 -7318 3020 -6942
rect 2962 -7330 3020 -7318
rect 3060 -6942 3118 -6930
rect 3060 -7318 3072 -6942
rect 3106 -7318 3118 -6942
rect 3060 -7330 3118 -7318
rect 3158 -6942 3216 -6930
rect 3158 -7318 3170 -6942
rect 3204 -7318 3216 -6942
rect 3158 -7330 3216 -7318
rect 3256 -6942 3314 -6930
rect 3256 -7318 3268 -6942
rect 3302 -7318 3314 -6942
rect 3256 -7330 3314 -7318
rect 3354 -6942 3412 -6930
rect 3354 -7318 3366 -6942
rect 3400 -7318 3412 -6942
rect 3354 -7330 3412 -7318
rect 3452 -6942 3510 -6930
rect 3452 -7318 3464 -6942
rect 3498 -7318 3510 -6942
rect 3452 -7330 3510 -7318
rect 3550 -6942 3608 -6930
rect 3550 -7318 3562 -6942
rect 3596 -7318 3608 -6942
rect 3550 -7330 3608 -7318
rect 3648 -6942 3706 -6930
rect 3648 -7318 3660 -6942
rect 3694 -7318 3706 -6942
rect 3648 -7330 3706 -7318
rect 3746 -6942 3804 -6930
rect 3746 -7318 3758 -6942
rect 3792 -7318 3804 -6942
rect 3746 -7330 3804 -7318
rect 3844 -6942 3902 -6930
rect 3844 -7318 3856 -6942
rect 3890 -7318 3902 -6942
rect 3844 -7330 3902 -7318
rect 3942 -6942 4000 -6930
rect 3942 -7318 3954 -6942
rect 3988 -7318 4000 -6942
rect 3942 -7330 4000 -7318
rect 1602 -8102 1664 -8090
rect 1602 -8478 1614 -8102
rect 1648 -8478 1664 -8102
rect 1602 -8490 1664 -8478
rect 1694 -8102 1760 -8090
rect 1694 -8478 1710 -8102
rect 1744 -8478 1760 -8102
rect 1694 -8490 1760 -8478
rect 1790 -8102 1856 -8090
rect 1790 -8478 1806 -8102
rect 1840 -8478 1856 -8102
rect 1790 -8490 1856 -8478
rect 1886 -8102 1952 -8090
rect 1886 -8478 1902 -8102
rect 1936 -8478 1952 -8102
rect 1886 -8490 1952 -8478
rect 1982 -8102 2048 -8090
rect 1982 -8478 1998 -8102
rect 2032 -8478 2048 -8102
rect 1982 -8490 2048 -8478
rect 2078 -8102 2144 -8090
rect 2078 -8478 2094 -8102
rect 2128 -8478 2144 -8102
rect 2078 -8490 2144 -8478
rect 2174 -8102 2240 -8090
rect 2174 -8478 2190 -8102
rect 2224 -8478 2240 -8102
rect 2174 -8490 2240 -8478
rect 2270 -8102 2336 -8090
rect 2270 -8478 2286 -8102
rect 2320 -8478 2336 -8102
rect 2270 -8490 2336 -8478
rect 2366 -8102 2432 -8090
rect 2366 -8478 2382 -8102
rect 2416 -8478 2432 -8102
rect 2366 -8490 2432 -8478
rect 2462 -8102 2528 -8090
rect 2462 -8478 2478 -8102
rect 2512 -8478 2528 -8102
rect 2462 -8490 2528 -8478
rect 2558 -8102 2624 -8090
rect 2558 -8478 2574 -8102
rect 2608 -8478 2624 -8102
rect 2558 -8490 2624 -8478
rect 2654 -8102 2720 -8090
rect 2654 -8478 2670 -8102
rect 2704 -8478 2720 -8102
rect 2654 -8490 2720 -8478
rect 2750 -8102 2812 -8090
rect 2750 -8478 2766 -8102
rect 2800 -8478 2812 -8102
rect 2750 -8490 2812 -8478
rect 3498 -8102 3560 -8090
rect 3498 -8478 3510 -8102
rect 3544 -8478 3560 -8102
rect 3498 -8490 3560 -8478
rect 3590 -8102 3656 -8090
rect 3590 -8478 3606 -8102
rect 3640 -8478 3656 -8102
rect 3590 -8490 3656 -8478
rect 3686 -8102 3752 -8090
rect 3686 -8478 3702 -8102
rect 3736 -8478 3752 -8102
rect 3686 -8490 3752 -8478
rect 3782 -8102 3848 -8090
rect 3782 -8478 3798 -8102
rect 3832 -8478 3848 -8102
rect 3782 -8490 3848 -8478
rect 3878 -8102 3944 -8090
rect 3878 -8478 3894 -8102
rect 3928 -8478 3944 -8102
rect 3878 -8490 3944 -8478
rect 3974 -8102 4040 -8090
rect 3974 -8478 3990 -8102
rect 4024 -8478 4040 -8102
rect 3974 -8490 4040 -8478
rect 4070 -8102 4136 -8090
rect 4070 -8478 4086 -8102
rect 4120 -8478 4136 -8102
rect 4070 -8490 4136 -8478
rect 4166 -8102 4232 -8090
rect 4166 -8478 4182 -8102
rect 4216 -8478 4232 -8102
rect 4166 -8490 4232 -8478
rect 4262 -8102 4328 -8090
rect 4262 -8478 4278 -8102
rect 4312 -8478 4328 -8102
rect 4262 -8490 4328 -8478
rect 4358 -8102 4424 -8090
rect 4358 -8478 4374 -8102
rect 4408 -8478 4424 -8102
rect 4358 -8490 4424 -8478
rect 4454 -8102 4520 -8090
rect 4454 -8478 4470 -8102
rect 4504 -8478 4520 -8102
rect 4454 -8490 4520 -8478
rect 4550 -8102 4616 -8090
rect 4550 -8478 4566 -8102
rect 4600 -8478 4616 -8102
rect 4550 -8490 4616 -8478
rect 4646 -8102 4708 -8090
rect 4646 -8478 4662 -8102
rect 4696 -8478 4708 -8102
rect 4646 -8490 4708 -8478
rect -1208 -8868 -1146 -8856
rect -1208 -9244 -1196 -8868
rect -1162 -9244 -1146 -8868
rect -1208 -9256 -1146 -9244
rect -1116 -8868 -1050 -8856
rect -1116 -9244 -1100 -8868
rect -1066 -9244 -1050 -8868
rect -1116 -9256 -1050 -9244
rect -1020 -8868 -954 -8856
rect -1020 -9244 -1004 -8868
rect -970 -9244 -954 -8868
rect -1020 -9256 -954 -9244
rect -924 -8868 -858 -8856
rect -924 -9244 -908 -8868
rect -874 -9244 -858 -8868
rect -924 -9256 -858 -9244
rect -828 -8868 -762 -8856
rect -828 -9244 -812 -8868
rect -778 -9244 -762 -8868
rect -828 -9256 -762 -9244
rect -732 -8868 -666 -8856
rect -732 -9244 -716 -8868
rect -682 -9244 -666 -8868
rect -732 -9256 -666 -9244
rect -636 -8868 -570 -8856
rect -636 -9244 -620 -8868
rect -586 -9244 -570 -8868
rect -636 -9256 -570 -9244
rect -540 -8868 -474 -8856
rect -540 -9244 -524 -8868
rect -490 -9244 -474 -8868
rect -540 -9256 -474 -9244
rect -444 -8868 -378 -8856
rect -444 -9244 -428 -8868
rect -394 -9244 -378 -8868
rect -444 -9256 -378 -9244
rect -348 -8868 -282 -8856
rect -348 -9244 -332 -8868
rect -298 -9244 -282 -8868
rect -348 -9256 -282 -9244
rect -252 -8868 -186 -8856
rect -252 -9244 -236 -8868
rect -202 -9244 -186 -8868
rect -252 -9256 -186 -9244
rect -156 -8868 -90 -8856
rect -156 -9244 -140 -8868
rect -106 -9244 -90 -8868
rect -156 -9256 -90 -9244
rect -60 -8868 6 -8856
rect -60 -9244 -44 -8868
rect -10 -9244 6 -8868
rect -60 -9256 6 -9244
rect 36 -8868 102 -8856
rect 36 -9244 52 -8868
rect 86 -9244 102 -8868
rect 36 -9256 102 -9244
rect 132 -8868 198 -8856
rect 132 -9244 148 -8868
rect 182 -9244 198 -8868
rect 132 -9256 198 -9244
rect 228 -8868 294 -8856
rect 228 -9244 244 -8868
rect 278 -9244 294 -8868
rect 228 -9256 294 -9244
rect 324 -8868 390 -8856
rect 324 -9244 340 -8868
rect 374 -9244 390 -8868
rect 324 -9256 390 -9244
rect 420 -8868 486 -8856
rect 420 -9244 436 -8868
rect 470 -9244 486 -8868
rect 420 -9256 486 -9244
rect 516 -8868 582 -8856
rect 516 -9244 532 -8868
rect 566 -9244 582 -8868
rect 516 -9256 582 -9244
rect 612 -8868 678 -8856
rect 612 -9244 628 -8868
rect 662 -9244 678 -8868
rect 612 -9256 678 -9244
rect 708 -8868 774 -8856
rect 708 -9244 724 -8868
rect 758 -9244 774 -8868
rect 708 -9256 774 -9244
rect 804 -8868 870 -8856
rect 804 -9244 820 -8868
rect 854 -9244 870 -8868
rect 804 -9256 870 -9244
rect 900 -8868 966 -8856
rect 900 -9244 916 -8868
rect 950 -9244 966 -8868
rect 900 -9256 966 -9244
rect 996 -8868 1062 -8856
rect 996 -9244 1012 -8868
rect 1046 -9244 1062 -8868
rect 996 -9256 1062 -9244
rect 1092 -8868 1158 -8856
rect 1092 -9244 1108 -8868
rect 1142 -9244 1158 -8868
rect 1092 -9256 1158 -9244
rect 1188 -8868 1250 -8856
rect 1188 -9244 1204 -8868
rect 1238 -9244 1250 -8868
rect 1188 -9256 1250 -9244
rect -1208 -9486 -1146 -9474
rect -1208 -9862 -1196 -9486
rect -1162 -9862 -1146 -9486
rect -1208 -9874 -1146 -9862
rect -1116 -9486 -1050 -9474
rect -1116 -9862 -1100 -9486
rect -1066 -9862 -1050 -9486
rect -1116 -9874 -1050 -9862
rect -1020 -9486 -954 -9474
rect -1020 -9862 -1004 -9486
rect -970 -9862 -954 -9486
rect -1020 -9874 -954 -9862
rect -924 -9486 -858 -9474
rect -924 -9862 -908 -9486
rect -874 -9862 -858 -9486
rect -924 -9874 -858 -9862
rect -828 -9486 -762 -9474
rect -828 -9862 -812 -9486
rect -778 -9862 -762 -9486
rect -828 -9874 -762 -9862
rect -732 -9486 -666 -9474
rect -732 -9862 -716 -9486
rect -682 -9862 -666 -9486
rect -732 -9874 -666 -9862
rect -636 -9486 -570 -9474
rect -636 -9862 -620 -9486
rect -586 -9862 -570 -9486
rect -636 -9874 -570 -9862
rect -540 -9486 -474 -9474
rect -540 -9862 -524 -9486
rect -490 -9862 -474 -9486
rect -540 -9874 -474 -9862
rect -444 -9486 -378 -9474
rect -444 -9862 -428 -9486
rect -394 -9862 -378 -9486
rect -444 -9874 -378 -9862
rect -348 -9486 -282 -9474
rect -348 -9862 -332 -9486
rect -298 -9862 -282 -9486
rect -348 -9874 -282 -9862
rect -252 -9486 -186 -9474
rect -252 -9862 -236 -9486
rect -202 -9862 -186 -9486
rect -252 -9874 -186 -9862
rect -156 -9486 -90 -9474
rect -156 -9862 -140 -9486
rect -106 -9862 -90 -9486
rect -156 -9874 -90 -9862
rect -60 -9486 6 -9474
rect -60 -9862 -44 -9486
rect -10 -9862 6 -9486
rect -60 -9874 6 -9862
rect 36 -9486 102 -9474
rect 36 -9862 52 -9486
rect 86 -9862 102 -9486
rect 36 -9874 102 -9862
rect 132 -9486 198 -9474
rect 132 -9862 148 -9486
rect 182 -9862 198 -9486
rect 132 -9874 198 -9862
rect 228 -9486 294 -9474
rect 228 -9862 244 -9486
rect 278 -9862 294 -9486
rect 228 -9874 294 -9862
rect 324 -9486 390 -9474
rect 324 -9862 340 -9486
rect 374 -9862 390 -9486
rect 324 -9874 390 -9862
rect 420 -9486 486 -9474
rect 420 -9862 436 -9486
rect 470 -9862 486 -9486
rect 420 -9874 486 -9862
rect 516 -9486 582 -9474
rect 516 -9862 532 -9486
rect 566 -9862 582 -9486
rect 516 -9874 582 -9862
rect 612 -9486 678 -9474
rect 612 -9862 628 -9486
rect 662 -9862 678 -9486
rect 612 -9874 678 -9862
rect 708 -9486 774 -9474
rect 708 -9862 724 -9486
rect 758 -9862 774 -9486
rect 708 -9874 774 -9862
rect 804 -9486 870 -9474
rect 804 -9862 820 -9486
rect 854 -9862 870 -9486
rect 804 -9874 870 -9862
rect 900 -9486 966 -9474
rect 900 -9862 916 -9486
rect 950 -9862 966 -9486
rect 900 -9874 966 -9862
rect 996 -9486 1062 -9474
rect 996 -9862 1012 -9486
rect 1046 -9862 1062 -9486
rect 996 -9874 1062 -9862
rect 1092 -9486 1158 -9474
rect 1092 -9862 1108 -9486
rect 1142 -9862 1158 -9486
rect 1092 -9874 1158 -9862
rect 1188 -9486 1250 -9474
rect 1188 -9862 1204 -9486
rect 1238 -9862 1250 -9486
rect 1188 -9874 1250 -9862
rect -1208 -10104 -1146 -10092
rect -1208 -10480 -1196 -10104
rect -1162 -10480 -1146 -10104
rect -1208 -10492 -1146 -10480
rect -1116 -10104 -1050 -10092
rect -1116 -10480 -1100 -10104
rect -1066 -10480 -1050 -10104
rect -1116 -10492 -1050 -10480
rect -1020 -10104 -954 -10092
rect -1020 -10480 -1004 -10104
rect -970 -10480 -954 -10104
rect -1020 -10492 -954 -10480
rect -924 -10104 -858 -10092
rect -924 -10480 -908 -10104
rect -874 -10480 -858 -10104
rect -924 -10492 -858 -10480
rect -828 -10104 -762 -10092
rect -828 -10480 -812 -10104
rect -778 -10480 -762 -10104
rect -828 -10492 -762 -10480
rect -732 -10104 -666 -10092
rect -732 -10480 -716 -10104
rect -682 -10480 -666 -10104
rect -732 -10492 -666 -10480
rect -636 -10104 -570 -10092
rect -636 -10480 -620 -10104
rect -586 -10480 -570 -10104
rect -636 -10492 -570 -10480
rect -540 -10104 -474 -10092
rect -540 -10480 -524 -10104
rect -490 -10480 -474 -10104
rect -540 -10492 -474 -10480
rect -444 -10104 -378 -10092
rect -444 -10480 -428 -10104
rect -394 -10480 -378 -10104
rect -444 -10492 -378 -10480
rect -348 -10104 -282 -10092
rect -348 -10480 -332 -10104
rect -298 -10480 -282 -10104
rect -348 -10492 -282 -10480
rect -252 -10104 -186 -10092
rect -252 -10480 -236 -10104
rect -202 -10480 -186 -10104
rect -252 -10492 -186 -10480
rect -156 -10104 -90 -10092
rect -156 -10480 -140 -10104
rect -106 -10480 -90 -10104
rect -156 -10492 -90 -10480
rect -60 -10104 6 -10092
rect -60 -10480 -44 -10104
rect -10 -10480 6 -10104
rect -60 -10492 6 -10480
rect 36 -10104 102 -10092
rect 36 -10480 52 -10104
rect 86 -10480 102 -10104
rect 36 -10492 102 -10480
rect 132 -10104 198 -10092
rect 132 -10480 148 -10104
rect 182 -10480 198 -10104
rect 132 -10492 198 -10480
rect 228 -10104 294 -10092
rect 228 -10480 244 -10104
rect 278 -10480 294 -10104
rect 228 -10492 294 -10480
rect 324 -10104 390 -10092
rect 324 -10480 340 -10104
rect 374 -10480 390 -10104
rect 324 -10492 390 -10480
rect 420 -10104 486 -10092
rect 420 -10480 436 -10104
rect 470 -10480 486 -10104
rect 420 -10492 486 -10480
rect 516 -10104 582 -10092
rect 516 -10480 532 -10104
rect 566 -10480 582 -10104
rect 516 -10492 582 -10480
rect 612 -10104 678 -10092
rect 612 -10480 628 -10104
rect 662 -10480 678 -10104
rect 612 -10492 678 -10480
rect 708 -10104 774 -10092
rect 708 -10480 724 -10104
rect 758 -10480 774 -10104
rect 708 -10492 774 -10480
rect 804 -10104 870 -10092
rect 804 -10480 820 -10104
rect 854 -10480 870 -10104
rect 804 -10492 870 -10480
rect 900 -10104 966 -10092
rect 900 -10480 916 -10104
rect 950 -10480 966 -10104
rect 900 -10492 966 -10480
rect 996 -10104 1062 -10092
rect 996 -10480 1012 -10104
rect 1046 -10480 1062 -10104
rect 996 -10492 1062 -10480
rect 1092 -10104 1158 -10092
rect 1092 -10480 1108 -10104
rect 1142 -10480 1158 -10104
rect 1092 -10492 1158 -10480
rect 1188 -10104 1250 -10092
rect 1188 -10480 1204 -10104
rect 1238 -10480 1250 -10104
rect 1188 -10492 1250 -10480
rect -1208 -10722 -1146 -10710
rect -1208 -11098 -1196 -10722
rect -1162 -11098 -1146 -10722
rect -1208 -11110 -1146 -11098
rect -1116 -10722 -1050 -10710
rect -1116 -11098 -1100 -10722
rect -1066 -11098 -1050 -10722
rect -1116 -11110 -1050 -11098
rect -1020 -10722 -954 -10710
rect -1020 -11098 -1004 -10722
rect -970 -11098 -954 -10722
rect -1020 -11110 -954 -11098
rect -924 -10722 -858 -10710
rect -924 -11098 -908 -10722
rect -874 -11098 -858 -10722
rect -924 -11110 -858 -11098
rect -828 -10722 -762 -10710
rect -828 -11098 -812 -10722
rect -778 -11098 -762 -10722
rect -828 -11110 -762 -11098
rect -732 -10722 -666 -10710
rect -732 -11098 -716 -10722
rect -682 -11098 -666 -10722
rect -732 -11110 -666 -11098
rect -636 -10722 -570 -10710
rect -636 -11098 -620 -10722
rect -586 -11098 -570 -10722
rect -636 -11110 -570 -11098
rect -540 -10722 -474 -10710
rect -540 -11098 -524 -10722
rect -490 -11098 -474 -10722
rect -540 -11110 -474 -11098
rect -444 -10722 -378 -10710
rect -444 -11098 -428 -10722
rect -394 -11098 -378 -10722
rect -444 -11110 -378 -11098
rect -348 -10722 -282 -10710
rect -348 -11098 -332 -10722
rect -298 -11098 -282 -10722
rect -348 -11110 -282 -11098
rect -252 -10722 -186 -10710
rect -252 -11098 -236 -10722
rect -202 -11098 -186 -10722
rect -252 -11110 -186 -11098
rect -156 -10722 -90 -10710
rect -156 -11098 -140 -10722
rect -106 -11098 -90 -10722
rect -156 -11110 -90 -11098
rect -60 -10722 6 -10710
rect -60 -11098 -44 -10722
rect -10 -11098 6 -10722
rect -60 -11110 6 -11098
rect 36 -10722 102 -10710
rect 36 -11098 52 -10722
rect 86 -11098 102 -10722
rect 36 -11110 102 -11098
rect 132 -10722 198 -10710
rect 132 -11098 148 -10722
rect 182 -11098 198 -10722
rect 132 -11110 198 -11098
rect 228 -10722 294 -10710
rect 228 -11098 244 -10722
rect 278 -11098 294 -10722
rect 228 -11110 294 -11098
rect 324 -10722 390 -10710
rect 324 -11098 340 -10722
rect 374 -11098 390 -10722
rect 324 -11110 390 -11098
rect 420 -10722 486 -10710
rect 420 -11098 436 -10722
rect 470 -11098 486 -10722
rect 420 -11110 486 -11098
rect 516 -10722 582 -10710
rect 516 -11098 532 -10722
rect 566 -11098 582 -10722
rect 516 -11110 582 -11098
rect 612 -10722 678 -10710
rect 612 -11098 628 -10722
rect 662 -11098 678 -10722
rect 612 -11110 678 -11098
rect 708 -10722 774 -10710
rect 708 -11098 724 -10722
rect 758 -11098 774 -10722
rect 708 -11110 774 -11098
rect 804 -10722 870 -10710
rect 804 -11098 820 -10722
rect 854 -11098 870 -10722
rect 804 -11110 870 -11098
rect 900 -10722 966 -10710
rect 900 -11098 916 -10722
rect 950 -11098 966 -10722
rect 900 -11110 966 -11098
rect 996 -10722 1062 -10710
rect 996 -11098 1012 -10722
rect 1046 -11098 1062 -10722
rect 996 -11110 1062 -11098
rect 1092 -10722 1158 -10710
rect 1092 -11098 1108 -10722
rect 1142 -11098 1158 -10722
rect 1092 -11110 1158 -11098
rect 1188 -10722 1250 -10710
rect 1188 -11098 1204 -10722
rect 1238 -11098 1250 -10722
rect 1188 -11110 1250 -11098
rect 1602 -8922 1660 -8910
rect 1602 -9298 1614 -8922
rect 1648 -9298 1660 -8922
rect 1602 -9310 1660 -9298
rect 1860 -8922 1918 -8910
rect 1860 -9298 1872 -8922
rect 1906 -9298 1918 -8922
rect 1860 -9310 1918 -9298
rect 2118 -8922 2176 -8910
rect 2118 -9298 2130 -8922
rect 2164 -9298 2176 -8922
rect 2118 -9310 2176 -9298
rect 2376 -8922 2434 -8910
rect 2376 -9298 2388 -8922
rect 2422 -9298 2434 -8922
rect 2376 -9310 2434 -9298
rect 2634 -8922 2692 -8910
rect 2634 -9298 2646 -8922
rect 2680 -9298 2692 -8922
rect 2634 -9310 2692 -9298
rect 2892 -8922 2950 -8910
rect 2892 -9298 2904 -8922
rect 2938 -9298 2950 -8922
rect 2892 -9310 2950 -9298
rect 3150 -8922 3208 -8910
rect 3150 -9298 3162 -8922
rect 3196 -9298 3208 -8922
rect 3150 -9310 3208 -9298
rect 3498 -8922 3556 -8910
rect 3498 -9298 3510 -8922
rect 3544 -9298 3556 -8922
rect 3498 -9310 3556 -9298
rect 3756 -8922 3814 -8910
rect 3756 -9298 3768 -8922
rect 3802 -9298 3814 -8922
rect 3756 -9310 3814 -9298
rect 4014 -8922 4072 -8910
rect 4014 -9298 4026 -8922
rect 4060 -9298 4072 -8922
rect 4014 -9310 4072 -9298
rect 4272 -8922 4330 -8910
rect 4272 -9298 4284 -8922
rect 4318 -9298 4330 -8922
rect 4272 -9310 4330 -9298
rect 4530 -8922 4588 -8910
rect 4530 -9298 4542 -8922
rect 4576 -9298 4588 -8922
rect 4530 -9310 4588 -9298
rect 4788 -8922 4846 -8910
rect 4788 -9298 4800 -8922
rect 4834 -9298 4846 -8922
rect 4788 -9310 4846 -9298
rect 5046 -8922 5104 -8910
rect 5046 -9298 5058 -8922
rect 5092 -9298 5104 -8922
rect 5046 -9310 5104 -9298
rect 5448 -8922 5510 -8910
rect 5448 -9298 5460 -8922
rect 5494 -9298 5510 -8922
rect 5448 -9310 5510 -9298
rect 5540 -8922 5606 -8910
rect 5540 -9298 5556 -8922
rect 5590 -9298 5606 -8922
rect 5540 -9310 5606 -9298
rect 5636 -8922 5702 -8910
rect 5636 -9298 5652 -8922
rect 5686 -9298 5702 -8922
rect 5636 -9310 5702 -9298
rect 5732 -8922 5798 -8910
rect 5732 -9298 5748 -8922
rect 5782 -9298 5798 -8922
rect 5732 -9310 5798 -9298
rect 5828 -8922 5894 -8910
rect 5828 -9298 5844 -8922
rect 5878 -9298 5894 -8922
rect 5828 -9310 5894 -9298
rect 5924 -8922 5986 -8910
rect 5924 -9298 5940 -8922
rect 5974 -9298 5986 -8922
rect 5924 -9310 5986 -9298
rect 6318 -10782 6376 -10770
rect 6318 -10858 6330 -10782
rect 6364 -10858 6376 -10782
rect 6318 -10870 6376 -10858
rect 6576 -10782 6634 -10770
rect 6576 -10858 6588 -10782
rect 6622 -10858 6634 -10782
rect 6576 -10870 6634 -10858
<< pdiff >>
rect -1188 2533 -1130 2545
rect -1188 2157 -1176 2533
rect -1142 2157 -1130 2533
rect -1188 2145 -1130 2157
rect -1090 2533 -1032 2545
rect -1090 2157 -1078 2533
rect -1044 2157 -1032 2533
rect -1090 2145 -1032 2157
rect -992 2533 -934 2545
rect -992 2157 -980 2533
rect -946 2157 -934 2533
rect -992 2145 -934 2157
rect -894 2533 -836 2545
rect -894 2157 -882 2533
rect -848 2157 -836 2533
rect -894 2145 -836 2157
rect -796 2533 -738 2545
rect -796 2157 -784 2533
rect -750 2157 -738 2533
rect -796 2145 -738 2157
rect -698 2533 -640 2545
rect -698 2157 -686 2533
rect -652 2157 -640 2533
rect -698 2145 -640 2157
rect -600 2533 -542 2545
rect -600 2157 -588 2533
rect -554 2157 -542 2533
rect -600 2145 -542 2157
rect -502 2533 -444 2545
rect -502 2157 -490 2533
rect -456 2157 -444 2533
rect -502 2145 -444 2157
rect -404 2533 -346 2545
rect -404 2157 -392 2533
rect -358 2157 -346 2533
rect -404 2145 -346 2157
rect -306 2533 -248 2545
rect -306 2157 -294 2533
rect -260 2157 -248 2533
rect -306 2145 -248 2157
rect -208 2533 -150 2545
rect -208 2157 -196 2533
rect -162 2157 -150 2533
rect -208 2145 -150 2157
rect -110 2533 -52 2545
rect -110 2157 -98 2533
rect -64 2157 -52 2533
rect -110 2145 -52 2157
rect -12 2533 46 2545
rect -12 2157 0 2533
rect 34 2157 46 2533
rect -12 2145 46 2157
rect 86 2533 144 2545
rect 86 2157 98 2533
rect 132 2157 144 2533
rect 86 2145 144 2157
rect 184 2533 242 2545
rect 184 2157 196 2533
rect 230 2157 242 2533
rect 184 2145 242 2157
rect 282 2533 340 2545
rect 282 2157 294 2533
rect 328 2157 340 2533
rect 282 2145 340 2157
rect -1188 1897 -1130 1909
rect -1188 1521 -1176 1897
rect -1142 1521 -1130 1897
rect -1188 1509 -1130 1521
rect -1090 1897 -1032 1909
rect -1090 1521 -1078 1897
rect -1044 1521 -1032 1897
rect -1090 1509 -1032 1521
rect -992 1897 -934 1909
rect -992 1521 -980 1897
rect -946 1521 -934 1897
rect -992 1509 -934 1521
rect -894 1897 -836 1909
rect -894 1521 -882 1897
rect -848 1521 -836 1897
rect -894 1509 -836 1521
rect -796 1897 -738 1909
rect -796 1521 -784 1897
rect -750 1521 -738 1897
rect -796 1509 -738 1521
rect -698 1897 -640 1909
rect -698 1521 -686 1897
rect -652 1521 -640 1897
rect -698 1509 -640 1521
rect -600 1897 -542 1909
rect -600 1521 -588 1897
rect -554 1521 -542 1897
rect -600 1509 -542 1521
rect -502 1897 -444 1909
rect -502 1521 -490 1897
rect -456 1521 -444 1897
rect -502 1509 -444 1521
rect -404 1897 -346 1909
rect -404 1521 -392 1897
rect -358 1521 -346 1897
rect -404 1509 -346 1521
rect -306 1897 -248 1909
rect -306 1521 -294 1897
rect -260 1521 -248 1897
rect -306 1509 -248 1521
rect -208 1897 -150 1909
rect -208 1521 -196 1897
rect -162 1521 -150 1897
rect -208 1509 -150 1521
rect -110 1897 -52 1909
rect -110 1521 -98 1897
rect -64 1521 -52 1897
rect -110 1509 -52 1521
rect -12 1897 46 1909
rect -12 1521 0 1897
rect 34 1521 46 1897
rect -12 1509 46 1521
rect 86 1897 144 1909
rect 86 1521 98 1897
rect 132 1521 144 1897
rect 86 1509 144 1521
rect 184 1897 242 1909
rect 184 1521 196 1897
rect 230 1521 242 1897
rect 184 1509 242 1521
rect 282 1897 340 1909
rect 282 1521 294 1897
rect 328 1521 340 1897
rect 282 1509 340 1521
rect 610 2533 668 2545
rect 610 2157 622 2533
rect 656 2157 668 2533
rect 610 2145 668 2157
rect 708 2533 766 2545
rect 708 2157 720 2533
rect 754 2157 766 2533
rect 708 2145 766 2157
rect 806 2533 864 2545
rect 806 2157 818 2533
rect 852 2157 864 2533
rect 806 2145 864 2157
rect 904 2533 962 2545
rect 904 2157 916 2533
rect 950 2157 962 2533
rect 904 2145 962 2157
rect 1002 2533 1060 2545
rect 1002 2157 1014 2533
rect 1048 2157 1060 2533
rect 1002 2145 1060 2157
rect 1100 2533 1158 2545
rect 1100 2157 1112 2533
rect 1146 2157 1158 2533
rect 1100 2145 1158 2157
rect 1198 2533 1256 2545
rect 1198 2157 1210 2533
rect 1244 2157 1256 2533
rect 1198 2145 1256 2157
rect 1296 2533 1354 2545
rect 1296 2157 1308 2533
rect 1342 2157 1354 2533
rect 1296 2145 1354 2157
rect 1394 2533 1452 2545
rect 1394 2157 1406 2533
rect 1440 2157 1452 2533
rect 1394 2145 1452 2157
rect 1492 2533 1550 2545
rect 1492 2157 1504 2533
rect 1538 2157 1550 2533
rect 1492 2145 1550 2157
rect 1590 2533 1648 2545
rect 1590 2157 1602 2533
rect 1636 2157 1648 2533
rect 1590 2145 1648 2157
rect 1688 2533 1746 2545
rect 1688 2157 1700 2533
rect 1734 2157 1746 2533
rect 1688 2145 1746 2157
rect 1786 2533 1844 2545
rect 1786 2157 1798 2533
rect 1832 2157 1844 2533
rect 1786 2145 1844 2157
rect 1884 2533 1942 2545
rect 1884 2157 1896 2533
rect 1930 2157 1942 2533
rect 1884 2145 1942 2157
rect 1982 2533 2040 2545
rect 1982 2157 1994 2533
rect 2028 2157 2040 2533
rect 1982 2145 2040 2157
rect 2080 2533 2138 2545
rect 2080 2157 2092 2533
rect 2126 2157 2138 2533
rect 2080 2145 2138 2157
rect 610 1897 668 1909
rect 610 1521 622 1897
rect 656 1521 668 1897
rect 610 1509 668 1521
rect 708 1897 766 1909
rect 708 1521 720 1897
rect 754 1521 766 1897
rect 708 1509 766 1521
rect 806 1897 864 1909
rect 806 1521 818 1897
rect 852 1521 864 1897
rect 806 1509 864 1521
rect 904 1897 962 1909
rect 904 1521 916 1897
rect 950 1521 962 1897
rect 904 1509 962 1521
rect 1002 1897 1060 1909
rect 1002 1521 1014 1897
rect 1048 1521 1060 1897
rect 1002 1509 1060 1521
rect 1100 1897 1158 1909
rect 1100 1521 1112 1897
rect 1146 1521 1158 1897
rect 1100 1509 1158 1521
rect 1198 1897 1256 1909
rect 1198 1521 1210 1897
rect 1244 1521 1256 1897
rect 1198 1509 1256 1521
rect 1296 1897 1354 1909
rect 1296 1521 1308 1897
rect 1342 1521 1354 1897
rect 1296 1509 1354 1521
rect 1394 1897 1452 1909
rect 1394 1521 1406 1897
rect 1440 1521 1452 1897
rect 1394 1509 1452 1521
rect 1492 1897 1550 1909
rect 1492 1521 1504 1897
rect 1538 1521 1550 1897
rect 1492 1509 1550 1521
rect 1590 1897 1648 1909
rect 1590 1521 1602 1897
rect 1636 1521 1648 1897
rect 1590 1509 1648 1521
rect 1688 1897 1746 1909
rect 1688 1521 1700 1897
rect 1734 1521 1746 1897
rect 1688 1509 1746 1521
rect 1786 1897 1844 1909
rect 1786 1521 1798 1897
rect 1832 1521 1844 1897
rect 1786 1509 1844 1521
rect 1884 1897 1942 1909
rect 1884 1521 1896 1897
rect 1930 1521 1942 1897
rect 1884 1509 1942 1521
rect 1982 1897 2040 1909
rect 1982 1521 1994 1897
rect 2028 1521 2040 1897
rect 1982 1509 2040 1521
rect 2080 1897 2138 1909
rect 2080 1521 2092 1897
rect 2126 1521 2138 1897
rect 2080 1509 2138 1521
rect 2412 1881 2470 1893
rect 2412 1505 2424 1881
rect 2458 1505 2470 1881
rect 2412 1493 2470 1505
rect 2570 1881 2628 1893
rect 2570 1505 2582 1881
rect 2616 1505 2628 1881
rect 2570 1493 2628 1505
rect 2728 1881 2786 1893
rect 2728 1505 2740 1881
rect 2774 1505 2786 1881
rect 2728 1493 2786 1505
rect 2886 1881 2944 1893
rect 2886 1505 2898 1881
rect 2932 1505 2944 1881
rect 2886 1493 2944 1505
rect 3044 1881 3102 1893
rect 3044 1505 3056 1881
rect 3090 1505 3102 1881
rect 3044 1493 3102 1505
rect 3202 1881 3260 1893
rect 3202 1505 3214 1881
rect 3248 1505 3260 1881
rect 3202 1493 3260 1505
rect 3360 1881 3418 1893
rect 3360 1505 3372 1881
rect 3406 1505 3418 1881
rect 3360 1493 3418 1505
rect 3518 1881 3576 1893
rect 3518 1505 3530 1881
rect 3564 1505 3576 1881
rect 3518 1493 3576 1505
rect 3676 1881 3734 1893
rect 3676 1505 3688 1881
rect 3722 1505 3734 1881
rect 3676 1493 3734 1505
rect 3834 1881 3892 1893
rect 3834 1505 3846 1881
rect 3880 1505 3892 1881
rect 3834 1493 3892 1505
rect 3992 1881 4050 1893
rect 3992 1505 4004 1881
rect 4038 1505 4050 1881
rect 3992 1493 4050 1505
rect -1188 -4537 -1130 -4525
rect -1188 -4913 -1176 -4537
rect -1142 -4913 -1130 -4537
rect -1188 -4925 -1130 -4913
rect -1090 -4537 -1032 -4525
rect -1090 -4913 -1078 -4537
rect -1044 -4913 -1032 -4537
rect -1090 -4925 -1032 -4913
rect -992 -4537 -934 -4525
rect -992 -4913 -980 -4537
rect -946 -4913 -934 -4537
rect -992 -4925 -934 -4913
rect -894 -4537 -836 -4525
rect -894 -4913 -882 -4537
rect -848 -4913 -836 -4537
rect -894 -4925 -836 -4913
rect -796 -4537 -738 -4525
rect -796 -4913 -784 -4537
rect -750 -4913 -738 -4537
rect -796 -4925 -738 -4913
rect -698 -4537 -640 -4525
rect -698 -4913 -686 -4537
rect -652 -4913 -640 -4537
rect -698 -4925 -640 -4913
rect -600 -4537 -542 -4525
rect -600 -4913 -588 -4537
rect -554 -4913 -542 -4537
rect -600 -4925 -542 -4913
rect -502 -4537 -444 -4525
rect -502 -4913 -490 -4537
rect -456 -4913 -444 -4537
rect -502 -4925 -444 -4913
rect -404 -4537 -346 -4525
rect -404 -4913 -392 -4537
rect -358 -4913 -346 -4537
rect -404 -4925 -346 -4913
rect -306 -4537 -248 -4525
rect -306 -4913 -294 -4537
rect -260 -4913 -248 -4537
rect -306 -4925 -248 -4913
rect -208 -4537 -150 -4525
rect -208 -4913 -196 -4537
rect -162 -4913 -150 -4537
rect -208 -4925 -150 -4913
rect -110 -4537 -52 -4525
rect -110 -4913 -98 -4537
rect -64 -4913 -52 -4537
rect -110 -4925 -52 -4913
rect -12 -4537 46 -4525
rect -12 -4913 0 -4537
rect 34 -4913 46 -4537
rect -12 -4925 46 -4913
rect 86 -4537 144 -4525
rect 86 -4913 98 -4537
rect 132 -4913 144 -4537
rect 86 -4925 144 -4913
rect 184 -4537 242 -4525
rect 184 -4913 196 -4537
rect 230 -4913 242 -4537
rect 184 -4925 242 -4913
rect 282 -4537 340 -4525
rect 282 -4913 294 -4537
rect 328 -4913 340 -4537
rect 282 -4925 340 -4913
rect -1188 -5173 -1130 -5161
rect -1188 -5549 -1176 -5173
rect -1142 -5549 -1130 -5173
rect -1188 -5561 -1130 -5549
rect -1090 -5173 -1032 -5161
rect -1090 -5549 -1078 -5173
rect -1044 -5549 -1032 -5173
rect -1090 -5561 -1032 -5549
rect -992 -5173 -934 -5161
rect -992 -5549 -980 -5173
rect -946 -5549 -934 -5173
rect -992 -5561 -934 -5549
rect -894 -5173 -836 -5161
rect -894 -5549 -882 -5173
rect -848 -5549 -836 -5173
rect -894 -5561 -836 -5549
rect -796 -5173 -738 -5161
rect -796 -5549 -784 -5173
rect -750 -5549 -738 -5173
rect -796 -5561 -738 -5549
rect -698 -5173 -640 -5161
rect -698 -5549 -686 -5173
rect -652 -5549 -640 -5173
rect -698 -5561 -640 -5549
rect -600 -5173 -542 -5161
rect -600 -5549 -588 -5173
rect -554 -5549 -542 -5173
rect -600 -5561 -542 -5549
rect -502 -5173 -444 -5161
rect -502 -5549 -490 -5173
rect -456 -5549 -444 -5173
rect -502 -5561 -444 -5549
rect -404 -5173 -346 -5161
rect -404 -5549 -392 -5173
rect -358 -5549 -346 -5173
rect -404 -5561 -346 -5549
rect -306 -5173 -248 -5161
rect -306 -5549 -294 -5173
rect -260 -5549 -248 -5173
rect -306 -5561 -248 -5549
rect -208 -5173 -150 -5161
rect -208 -5549 -196 -5173
rect -162 -5549 -150 -5173
rect -208 -5561 -150 -5549
rect -110 -5173 -52 -5161
rect -110 -5549 -98 -5173
rect -64 -5549 -52 -5173
rect -110 -5561 -52 -5549
rect -12 -5173 46 -5161
rect -12 -5549 0 -5173
rect 34 -5549 46 -5173
rect -12 -5561 46 -5549
rect 86 -5173 144 -5161
rect 86 -5549 98 -5173
rect 132 -5549 144 -5173
rect 86 -5561 144 -5549
rect 184 -5173 242 -5161
rect 184 -5549 196 -5173
rect 230 -5549 242 -5173
rect 184 -5561 242 -5549
rect 282 -5173 340 -5161
rect 282 -5549 294 -5173
rect 328 -5549 340 -5173
rect 282 -5561 340 -5549
rect 610 -4537 668 -4525
rect 610 -4913 622 -4537
rect 656 -4913 668 -4537
rect 610 -4925 668 -4913
rect 708 -4537 766 -4525
rect 708 -4913 720 -4537
rect 754 -4913 766 -4537
rect 708 -4925 766 -4913
rect 806 -4537 864 -4525
rect 806 -4913 818 -4537
rect 852 -4913 864 -4537
rect 806 -4925 864 -4913
rect 904 -4537 962 -4525
rect 904 -4913 916 -4537
rect 950 -4913 962 -4537
rect 904 -4925 962 -4913
rect 1002 -4537 1060 -4525
rect 1002 -4913 1014 -4537
rect 1048 -4913 1060 -4537
rect 1002 -4925 1060 -4913
rect 1100 -4537 1158 -4525
rect 1100 -4913 1112 -4537
rect 1146 -4913 1158 -4537
rect 1100 -4925 1158 -4913
rect 1198 -4537 1256 -4525
rect 1198 -4913 1210 -4537
rect 1244 -4913 1256 -4537
rect 1198 -4925 1256 -4913
rect 1296 -4537 1354 -4525
rect 1296 -4913 1308 -4537
rect 1342 -4913 1354 -4537
rect 1296 -4925 1354 -4913
rect 1394 -4537 1452 -4525
rect 1394 -4913 1406 -4537
rect 1440 -4913 1452 -4537
rect 1394 -4925 1452 -4913
rect 1492 -4537 1550 -4525
rect 1492 -4913 1504 -4537
rect 1538 -4913 1550 -4537
rect 1492 -4925 1550 -4913
rect 1590 -4537 1648 -4525
rect 1590 -4913 1602 -4537
rect 1636 -4913 1648 -4537
rect 1590 -4925 1648 -4913
rect 1688 -4537 1746 -4525
rect 1688 -4913 1700 -4537
rect 1734 -4913 1746 -4537
rect 1688 -4925 1746 -4913
rect 1786 -4537 1844 -4525
rect 1786 -4913 1798 -4537
rect 1832 -4913 1844 -4537
rect 1786 -4925 1844 -4913
rect 1884 -4537 1942 -4525
rect 1884 -4913 1896 -4537
rect 1930 -4913 1942 -4537
rect 1884 -4925 1942 -4913
rect 1982 -4537 2040 -4525
rect 1982 -4913 1994 -4537
rect 2028 -4913 2040 -4537
rect 1982 -4925 2040 -4913
rect 2080 -4537 2138 -4525
rect 2080 -4913 2092 -4537
rect 2126 -4913 2138 -4537
rect 2080 -4925 2138 -4913
rect 610 -5173 668 -5161
rect 610 -5549 622 -5173
rect 656 -5549 668 -5173
rect 610 -5561 668 -5549
rect 708 -5173 766 -5161
rect 708 -5549 720 -5173
rect 754 -5549 766 -5173
rect 708 -5561 766 -5549
rect 806 -5173 864 -5161
rect 806 -5549 818 -5173
rect 852 -5549 864 -5173
rect 806 -5561 864 -5549
rect 904 -5173 962 -5161
rect 904 -5549 916 -5173
rect 950 -5549 962 -5173
rect 904 -5561 962 -5549
rect 1002 -5173 1060 -5161
rect 1002 -5549 1014 -5173
rect 1048 -5549 1060 -5173
rect 1002 -5561 1060 -5549
rect 1100 -5173 1158 -5161
rect 1100 -5549 1112 -5173
rect 1146 -5549 1158 -5173
rect 1100 -5561 1158 -5549
rect 1198 -5173 1256 -5161
rect 1198 -5549 1210 -5173
rect 1244 -5549 1256 -5173
rect 1198 -5561 1256 -5549
rect 1296 -5173 1354 -5161
rect 1296 -5549 1308 -5173
rect 1342 -5549 1354 -5173
rect 1296 -5561 1354 -5549
rect 1394 -5173 1452 -5161
rect 1394 -5549 1406 -5173
rect 1440 -5549 1452 -5173
rect 1394 -5561 1452 -5549
rect 1492 -5173 1550 -5161
rect 1492 -5549 1504 -5173
rect 1538 -5549 1550 -5173
rect 1492 -5561 1550 -5549
rect 1590 -5173 1648 -5161
rect 1590 -5549 1602 -5173
rect 1636 -5549 1648 -5173
rect 1590 -5561 1648 -5549
rect 1688 -5173 1746 -5161
rect 1688 -5549 1700 -5173
rect 1734 -5549 1746 -5173
rect 1688 -5561 1746 -5549
rect 1786 -5173 1844 -5161
rect 1786 -5549 1798 -5173
rect 1832 -5549 1844 -5173
rect 1786 -5561 1844 -5549
rect 1884 -5173 1942 -5161
rect 1884 -5549 1896 -5173
rect 1930 -5549 1942 -5173
rect 1884 -5561 1942 -5549
rect 1982 -5173 2040 -5161
rect 1982 -5549 1994 -5173
rect 2028 -5549 2040 -5173
rect 1982 -5561 2040 -5549
rect 2080 -5173 2138 -5161
rect 2080 -5549 2092 -5173
rect 2126 -5549 2138 -5173
rect 2080 -5561 2138 -5549
rect 2412 -5189 2470 -5177
rect 2412 -5565 2424 -5189
rect 2458 -5565 2470 -5189
rect 2412 -5577 2470 -5565
rect 2570 -5189 2628 -5177
rect 2570 -5565 2582 -5189
rect 2616 -5565 2628 -5189
rect 2570 -5577 2628 -5565
rect 2728 -5189 2786 -5177
rect 2728 -5565 2740 -5189
rect 2774 -5565 2786 -5189
rect 2728 -5577 2786 -5565
rect 2886 -5189 2944 -5177
rect 2886 -5565 2898 -5189
rect 2932 -5565 2944 -5189
rect 2886 -5577 2944 -5565
rect 3044 -5189 3102 -5177
rect 3044 -5565 3056 -5189
rect 3090 -5565 3102 -5189
rect 3044 -5577 3102 -5565
rect 3202 -5189 3260 -5177
rect 3202 -5565 3214 -5189
rect 3248 -5565 3260 -5189
rect 3202 -5577 3260 -5565
rect 3360 -5189 3418 -5177
rect 3360 -5565 3372 -5189
rect 3406 -5565 3418 -5189
rect 3360 -5577 3418 -5565
rect 3518 -5189 3576 -5177
rect 3518 -5565 3530 -5189
rect 3564 -5565 3576 -5189
rect 3518 -5577 3576 -5565
rect 3676 -5189 3734 -5177
rect 3676 -5565 3688 -5189
rect 3722 -5565 3734 -5189
rect 3676 -5577 3734 -5565
rect 3834 -5189 3892 -5177
rect 3834 -5565 3846 -5189
rect 3880 -5565 3892 -5189
rect 3834 -5577 3892 -5565
rect 3992 -5189 4050 -5177
rect 3992 -5565 4004 -5189
rect 4038 -5565 4050 -5189
rect 3992 -5577 4050 -5565
rect 6318 -10223 6376 -10211
rect 6318 -10299 6330 -10223
rect 6364 -10299 6376 -10223
rect 6318 -10311 6376 -10299
rect 6576 -10223 6634 -10211
rect 6576 -10299 6588 -10223
rect 6622 -10299 6634 -10223
rect 6576 -10311 6634 -10299
<< ndiffc >>
rect -1176 690 -1142 1066
rect -1078 690 -1044 1066
rect -980 690 -946 1066
rect -882 690 -848 1066
rect -784 690 -750 1066
rect -686 690 -652 1066
rect -588 690 -554 1066
rect -490 690 -456 1066
rect -392 690 -358 1066
rect -294 690 -260 1066
rect -196 690 -162 1066
rect -98 690 -64 1066
rect 0 690 34 1066
rect 98 690 132 1066
rect 196 690 230 1066
rect 294 690 328 1066
rect 392 690 426 1066
rect 490 690 524 1066
rect 588 690 622 1066
rect 686 690 720 1066
rect 784 690 818 1066
rect 882 690 916 1066
rect 980 690 1014 1066
rect 1078 690 1112 1066
rect 1176 690 1210 1066
rect 1274 690 1308 1066
rect -1176 72 -1142 448
rect -1078 72 -1044 448
rect -980 72 -946 448
rect -882 72 -848 448
rect -784 72 -750 448
rect -686 72 -652 448
rect -588 72 -554 448
rect -490 72 -456 448
rect -392 72 -358 448
rect -294 72 -260 448
rect -196 72 -162 448
rect -98 72 -64 448
rect 0 72 34 448
rect 98 72 132 448
rect 196 72 230 448
rect 294 72 328 448
rect 392 72 426 448
rect 490 72 524 448
rect 588 72 622 448
rect 686 72 720 448
rect 784 72 818 448
rect 882 72 916 448
rect 980 72 1014 448
rect 1078 72 1112 448
rect 1176 72 1210 448
rect 1274 72 1308 448
rect -1176 -754 -1142 -378
rect -1078 -754 -1044 -378
rect -980 -754 -946 -378
rect -882 -754 -848 -378
rect -784 -754 -750 -378
rect -686 -754 -652 -378
rect -588 -754 -554 -378
rect -490 -754 -456 -378
rect -392 -754 -358 -378
rect -294 -754 -260 -378
rect -196 -754 -162 -378
rect -98 -754 -64 -378
rect 0 -754 34 -378
rect 98 -754 132 -378
rect 196 -754 230 -378
rect 294 -754 328 -378
rect 392 -754 426 -378
rect 490 -754 524 -378
rect 588 -754 622 -378
rect 686 -754 720 -378
rect 784 -754 818 -378
rect 882 -754 916 -378
rect 980 -754 1014 -378
rect 1078 -754 1112 -378
rect 1176 -754 1210 -378
rect 1274 -754 1308 -378
rect -1176 -1372 -1142 -996
rect -1078 -1372 -1044 -996
rect -980 -1372 -946 -996
rect -882 -1372 -848 -996
rect -784 -1372 -750 -996
rect -686 -1372 -652 -996
rect -588 -1372 -554 -996
rect -490 -1372 -456 -996
rect -392 -1372 -358 -996
rect -294 -1372 -260 -996
rect -196 -1372 -162 -996
rect -98 -1372 -64 -996
rect 0 -1372 34 -996
rect 98 -1372 132 -996
rect 196 -1372 230 -996
rect 294 -1372 328 -996
rect 392 -1372 426 -996
rect 490 -1372 524 -996
rect 588 -1372 622 -996
rect 686 -1372 720 -996
rect 784 -1372 818 -996
rect 882 -1372 916 -996
rect 980 -1372 1014 -996
rect 1078 -1372 1112 -996
rect 1176 -1372 1210 -996
rect 1274 -1372 1308 -996
rect 2484 370 2518 746
rect 2582 370 2616 746
rect 2680 370 2714 746
rect 2778 370 2812 746
rect 2876 370 2910 746
rect 2974 370 3008 746
rect 3072 370 3106 746
rect 3170 370 3204 746
rect 3268 370 3302 746
rect 3366 370 3400 746
rect 3464 370 3498 746
rect 3562 370 3596 746
rect 3660 370 3694 746
rect 3758 370 3792 746
rect 3856 370 3890 746
rect 3954 370 3988 746
rect 2484 -248 2518 128
rect 2582 -248 2616 128
rect 2680 -248 2714 128
rect 2778 -248 2812 128
rect 2876 -248 2910 128
rect 2974 -248 3008 128
rect 3072 -248 3106 128
rect 3170 -248 3204 128
rect 3268 -248 3302 128
rect 3366 -248 3400 128
rect 3464 -248 3498 128
rect 3562 -248 3596 128
rect 3660 -248 3694 128
rect 3758 -248 3792 128
rect 3856 -248 3890 128
rect 3954 -248 3988 128
rect 1614 -1408 1648 -1032
rect 1710 -1408 1744 -1032
rect 1806 -1408 1840 -1032
rect 1902 -1408 1936 -1032
rect 1998 -1408 2032 -1032
rect 2094 -1408 2128 -1032
rect 2190 -1408 2224 -1032
rect 2286 -1408 2320 -1032
rect 2382 -1408 2416 -1032
rect 2478 -1408 2512 -1032
rect 2574 -1408 2608 -1032
rect 2670 -1408 2704 -1032
rect 2766 -1408 2800 -1032
rect -1196 -2174 -1162 -1798
rect -1100 -2174 -1066 -1798
rect -1004 -2174 -970 -1798
rect -908 -2174 -874 -1798
rect -812 -2174 -778 -1798
rect -716 -2174 -682 -1798
rect -620 -2174 -586 -1798
rect -524 -2174 -490 -1798
rect -428 -2174 -394 -1798
rect -332 -2174 -298 -1798
rect -236 -2174 -202 -1798
rect -140 -2174 -106 -1798
rect -44 -2174 -10 -1798
rect 52 -2174 86 -1798
rect 148 -2174 182 -1798
rect 244 -2174 278 -1798
rect 340 -2174 374 -1798
rect 436 -2174 470 -1798
rect 532 -2174 566 -1798
rect 628 -2174 662 -1798
rect 724 -2174 758 -1798
rect 820 -2174 854 -1798
rect 916 -2174 950 -1798
rect 1012 -2174 1046 -1798
rect 1108 -2174 1142 -1798
rect 1204 -2174 1238 -1798
rect -1196 -2792 -1162 -2416
rect -1100 -2792 -1066 -2416
rect -1004 -2792 -970 -2416
rect -908 -2792 -874 -2416
rect -812 -2792 -778 -2416
rect -716 -2792 -682 -2416
rect -620 -2792 -586 -2416
rect -524 -2792 -490 -2416
rect -428 -2792 -394 -2416
rect -332 -2792 -298 -2416
rect -236 -2792 -202 -2416
rect -140 -2792 -106 -2416
rect -44 -2792 -10 -2416
rect 52 -2792 86 -2416
rect 148 -2792 182 -2416
rect 244 -2792 278 -2416
rect 340 -2792 374 -2416
rect 436 -2792 470 -2416
rect 532 -2792 566 -2416
rect 628 -2792 662 -2416
rect 724 -2792 758 -2416
rect 820 -2792 854 -2416
rect 916 -2792 950 -2416
rect 1012 -2792 1046 -2416
rect 1108 -2792 1142 -2416
rect 1204 -2792 1238 -2416
rect -1196 -3410 -1162 -3034
rect -1100 -3410 -1066 -3034
rect -1004 -3410 -970 -3034
rect -908 -3410 -874 -3034
rect -812 -3410 -778 -3034
rect -716 -3410 -682 -3034
rect -620 -3410 -586 -3034
rect -524 -3410 -490 -3034
rect -428 -3410 -394 -3034
rect -332 -3410 -298 -3034
rect -236 -3410 -202 -3034
rect -140 -3410 -106 -3034
rect -44 -3410 -10 -3034
rect 52 -3410 86 -3034
rect 148 -3410 182 -3034
rect 244 -3410 278 -3034
rect 340 -3410 374 -3034
rect 436 -3410 470 -3034
rect 532 -3410 566 -3034
rect 628 -3410 662 -3034
rect 724 -3410 758 -3034
rect 820 -3410 854 -3034
rect 916 -3410 950 -3034
rect 1012 -3410 1046 -3034
rect 1108 -3410 1142 -3034
rect 1204 -3410 1238 -3034
rect -1196 -4028 -1162 -3652
rect -1100 -4028 -1066 -3652
rect -1004 -4028 -970 -3652
rect -908 -4028 -874 -3652
rect -812 -4028 -778 -3652
rect -716 -4028 -682 -3652
rect -620 -4028 -586 -3652
rect -524 -4028 -490 -3652
rect -428 -4028 -394 -3652
rect -332 -4028 -298 -3652
rect -236 -4028 -202 -3652
rect -140 -4028 -106 -3652
rect -44 -4028 -10 -3652
rect 52 -4028 86 -3652
rect 148 -4028 182 -3652
rect 244 -4028 278 -3652
rect 340 -4028 374 -3652
rect 436 -4028 470 -3652
rect 532 -4028 566 -3652
rect 628 -4028 662 -3652
rect 724 -4028 758 -3652
rect 820 -4028 854 -3652
rect 916 -4028 950 -3652
rect 1012 -4028 1046 -3652
rect 1108 -4028 1142 -3652
rect 1204 -4028 1238 -3652
rect 1614 -2228 1648 -1852
rect 1872 -2228 1906 -1852
rect 2130 -2228 2164 -1852
rect 2388 -2228 2422 -1852
rect 2646 -2228 2680 -1852
rect 2904 -2228 2938 -1852
rect 3162 -2228 3196 -1852
rect -1176 -6380 -1142 -6004
rect -1078 -6380 -1044 -6004
rect -980 -6380 -946 -6004
rect -882 -6380 -848 -6004
rect -784 -6380 -750 -6004
rect -686 -6380 -652 -6004
rect -588 -6380 -554 -6004
rect -490 -6380 -456 -6004
rect -392 -6380 -358 -6004
rect -294 -6380 -260 -6004
rect -196 -6380 -162 -6004
rect -98 -6380 -64 -6004
rect 0 -6380 34 -6004
rect 98 -6380 132 -6004
rect 196 -6380 230 -6004
rect 294 -6380 328 -6004
rect 392 -6380 426 -6004
rect 490 -6380 524 -6004
rect 588 -6380 622 -6004
rect 686 -6380 720 -6004
rect 784 -6380 818 -6004
rect 882 -6380 916 -6004
rect 980 -6380 1014 -6004
rect 1078 -6380 1112 -6004
rect 1176 -6380 1210 -6004
rect 1274 -6380 1308 -6004
rect -1176 -6998 -1142 -6622
rect -1078 -6998 -1044 -6622
rect -980 -6998 -946 -6622
rect -882 -6998 -848 -6622
rect -784 -6998 -750 -6622
rect -686 -6998 -652 -6622
rect -588 -6998 -554 -6622
rect -490 -6998 -456 -6622
rect -392 -6998 -358 -6622
rect -294 -6998 -260 -6622
rect -196 -6998 -162 -6622
rect -98 -6998 -64 -6622
rect 0 -6998 34 -6622
rect 98 -6998 132 -6622
rect 196 -6998 230 -6622
rect 294 -6998 328 -6622
rect 392 -6998 426 -6622
rect 490 -6998 524 -6622
rect 588 -6998 622 -6622
rect 686 -6998 720 -6622
rect 784 -6998 818 -6622
rect 882 -6998 916 -6622
rect 980 -6998 1014 -6622
rect 1078 -6998 1112 -6622
rect 1176 -6998 1210 -6622
rect 1274 -6998 1308 -6622
rect -1176 -7824 -1142 -7448
rect -1078 -7824 -1044 -7448
rect -980 -7824 -946 -7448
rect -882 -7824 -848 -7448
rect -784 -7824 -750 -7448
rect -686 -7824 -652 -7448
rect -588 -7824 -554 -7448
rect -490 -7824 -456 -7448
rect -392 -7824 -358 -7448
rect -294 -7824 -260 -7448
rect -196 -7824 -162 -7448
rect -98 -7824 -64 -7448
rect 0 -7824 34 -7448
rect 98 -7824 132 -7448
rect 196 -7824 230 -7448
rect 294 -7824 328 -7448
rect 392 -7824 426 -7448
rect 490 -7824 524 -7448
rect 588 -7824 622 -7448
rect 686 -7824 720 -7448
rect 784 -7824 818 -7448
rect 882 -7824 916 -7448
rect 980 -7824 1014 -7448
rect 1078 -7824 1112 -7448
rect 1176 -7824 1210 -7448
rect 1274 -7824 1308 -7448
rect -1176 -8442 -1142 -8066
rect -1078 -8442 -1044 -8066
rect -980 -8442 -946 -8066
rect -882 -8442 -848 -8066
rect -784 -8442 -750 -8066
rect -686 -8442 -652 -8066
rect -588 -8442 -554 -8066
rect -490 -8442 -456 -8066
rect -392 -8442 -358 -8066
rect -294 -8442 -260 -8066
rect -196 -8442 -162 -8066
rect -98 -8442 -64 -8066
rect 0 -8442 34 -8066
rect 98 -8442 132 -8066
rect 196 -8442 230 -8066
rect 294 -8442 328 -8066
rect 392 -8442 426 -8066
rect 490 -8442 524 -8066
rect 588 -8442 622 -8066
rect 686 -8442 720 -8066
rect 784 -8442 818 -8066
rect 882 -8442 916 -8066
rect 980 -8442 1014 -8066
rect 1078 -8442 1112 -8066
rect 1176 -8442 1210 -8066
rect 1274 -8442 1308 -8066
rect 2484 -6700 2518 -6324
rect 2582 -6700 2616 -6324
rect 2680 -6700 2714 -6324
rect 2778 -6700 2812 -6324
rect 2876 -6700 2910 -6324
rect 2974 -6700 3008 -6324
rect 3072 -6700 3106 -6324
rect 3170 -6700 3204 -6324
rect 3268 -6700 3302 -6324
rect 3366 -6700 3400 -6324
rect 3464 -6700 3498 -6324
rect 3562 -6700 3596 -6324
rect 3660 -6700 3694 -6324
rect 3758 -6700 3792 -6324
rect 3856 -6700 3890 -6324
rect 3954 -6700 3988 -6324
rect 2484 -7318 2518 -6942
rect 2582 -7318 2616 -6942
rect 2680 -7318 2714 -6942
rect 2778 -7318 2812 -6942
rect 2876 -7318 2910 -6942
rect 2974 -7318 3008 -6942
rect 3072 -7318 3106 -6942
rect 3170 -7318 3204 -6942
rect 3268 -7318 3302 -6942
rect 3366 -7318 3400 -6942
rect 3464 -7318 3498 -6942
rect 3562 -7318 3596 -6942
rect 3660 -7318 3694 -6942
rect 3758 -7318 3792 -6942
rect 3856 -7318 3890 -6942
rect 3954 -7318 3988 -6942
rect 1614 -8478 1648 -8102
rect 1710 -8478 1744 -8102
rect 1806 -8478 1840 -8102
rect 1902 -8478 1936 -8102
rect 1998 -8478 2032 -8102
rect 2094 -8478 2128 -8102
rect 2190 -8478 2224 -8102
rect 2286 -8478 2320 -8102
rect 2382 -8478 2416 -8102
rect 2478 -8478 2512 -8102
rect 2574 -8478 2608 -8102
rect 2670 -8478 2704 -8102
rect 2766 -8478 2800 -8102
rect 3510 -8478 3544 -8102
rect 3606 -8478 3640 -8102
rect 3702 -8478 3736 -8102
rect 3798 -8478 3832 -8102
rect 3894 -8478 3928 -8102
rect 3990 -8478 4024 -8102
rect 4086 -8478 4120 -8102
rect 4182 -8478 4216 -8102
rect 4278 -8478 4312 -8102
rect 4374 -8478 4408 -8102
rect 4470 -8478 4504 -8102
rect 4566 -8478 4600 -8102
rect 4662 -8478 4696 -8102
rect -1196 -9244 -1162 -8868
rect -1100 -9244 -1066 -8868
rect -1004 -9244 -970 -8868
rect -908 -9244 -874 -8868
rect -812 -9244 -778 -8868
rect -716 -9244 -682 -8868
rect -620 -9244 -586 -8868
rect -524 -9244 -490 -8868
rect -428 -9244 -394 -8868
rect -332 -9244 -298 -8868
rect -236 -9244 -202 -8868
rect -140 -9244 -106 -8868
rect -44 -9244 -10 -8868
rect 52 -9244 86 -8868
rect 148 -9244 182 -8868
rect 244 -9244 278 -8868
rect 340 -9244 374 -8868
rect 436 -9244 470 -8868
rect 532 -9244 566 -8868
rect 628 -9244 662 -8868
rect 724 -9244 758 -8868
rect 820 -9244 854 -8868
rect 916 -9244 950 -8868
rect 1012 -9244 1046 -8868
rect 1108 -9244 1142 -8868
rect 1204 -9244 1238 -8868
rect -1196 -9862 -1162 -9486
rect -1100 -9862 -1066 -9486
rect -1004 -9862 -970 -9486
rect -908 -9862 -874 -9486
rect -812 -9862 -778 -9486
rect -716 -9862 -682 -9486
rect -620 -9862 -586 -9486
rect -524 -9862 -490 -9486
rect -428 -9862 -394 -9486
rect -332 -9862 -298 -9486
rect -236 -9862 -202 -9486
rect -140 -9862 -106 -9486
rect -44 -9862 -10 -9486
rect 52 -9862 86 -9486
rect 148 -9862 182 -9486
rect 244 -9862 278 -9486
rect 340 -9862 374 -9486
rect 436 -9862 470 -9486
rect 532 -9862 566 -9486
rect 628 -9862 662 -9486
rect 724 -9862 758 -9486
rect 820 -9862 854 -9486
rect 916 -9862 950 -9486
rect 1012 -9862 1046 -9486
rect 1108 -9862 1142 -9486
rect 1204 -9862 1238 -9486
rect -1196 -10480 -1162 -10104
rect -1100 -10480 -1066 -10104
rect -1004 -10480 -970 -10104
rect -908 -10480 -874 -10104
rect -812 -10480 -778 -10104
rect -716 -10480 -682 -10104
rect -620 -10480 -586 -10104
rect -524 -10480 -490 -10104
rect -428 -10480 -394 -10104
rect -332 -10480 -298 -10104
rect -236 -10480 -202 -10104
rect -140 -10480 -106 -10104
rect -44 -10480 -10 -10104
rect 52 -10480 86 -10104
rect 148 -10480 182 -10104
rect 244 -10480 278 -10104
rect 340 -10480 374 -10104
rect 436 -10480 470 -10104
rect 532 -10480 566 -10104
rect 628 -10480 662 -10104
rect 724 -10480 758 -10104
rect 820 -10480 854 -10104
rect 916 -10480 950 -10104
rect 1012 -10480 1046 -10104
rect 1108 -10480 1142 -10104
rect 1204 -10480 1238 -10104
rect -1196 -11098 -1162 -10722
rect -1100 -11098 -1066 -10722
rect -1004 -11098 -970 -10722
rect -908 -11098 -874 -10722
rect -812 -11098 -778 -10722
rect -716 -11098 -682 -10722
rect -620 -11098 -586 -10722
rect -524 -11098 -490 -10722
rect -428 -11098 -394 -10722
rect -332 -11098 -298 -10722
rect -236 -11098 -202 -10722
rect -140 -11098 -106 -10722
rect -44 -11098 -10 -10722
rect 52 -11098 86 -10722
rect 148 -11098 182 -10722
rect 244 -11098 278 -10722
rect 340 -11098 374 -10722
rect 436 -11098 470 -10722
rect 532 -11098 566 -10722
rect 628 -11098 662 -10722
rect 724 -11098 758 -10722
rect 820 -11098 854 -10722
rect 916 -11098 950 -10722
rect 1012 -11098 1046 -10722
rect 1108 -11098 1142 -10722
rect 1204 -11098 1238 -10722
rect 1614 -9298 1648 -8922
rect 1872 -9298 1906 -8922
rect 2130 -9298 2164 -8922
rect 2388 -9298 2422 -8922
rect 2646 -9298 2680 -8922
rect 2904 -9298 2938 -8922
rect 3162 -9298 3196 -8922
rect 3510 -9298 3544 -8922
rect 3768 -9298 3802 -8922
rect 4026 -9298 4060 -8922
rect 4284 -9298 4318 -8922
rect 4542 -9298 4576 -8922
rect 4800 -9298 4834 -8922
rect 5058 -9298 5092 -8922
rect 5460 -9298 5494 -8922
rect 5556 -9298 5590 -8922
rect 5652 -9298 5686 -8922
rect 5748 -9298 5782 -8922
rect 5844 -9298 5878 -8922
rect 5940 -9298 5974 -8922
rect 6330 -10858 6364 -10782
rect 6588 -10858 6622 -10782
<< pdiffc >>
rect -1176 2157 -1142 2533
rect -1078 2157 -1044 2533
rect -980 2157 -946 2533
rect -882 2157 -848 2533
rect -784 2157 -750 2533
rect -686 2157 -652 2533
rect -588 2157 -554 2533
rect -490 2157 -456 2533
rect -392 2157 -358 2533
rect -294 2157 -260 2533
rect -196 2157 -162 2533
rect -98 2157 -64 2533
rect 0 2157 34 2533
rect 98 2157 132 2533
rect 196 2157 230 2533
rect 294 2157 328 2533
rect -1176 1521 -1142 1897
rect -1078 1521 -1044 1897
rect -980 1521 -946 1897
rect -882 1521 -848 1897
rect -784 1521 -750 1897
rect -686 1521 -652 1897
rect -588 1521 -554 1897
rect -490 1521 -456 1897
rect -392 1521 -358 1897
rect -294 1521 -260 1897
rect -196 1521 -162 1897
rect -98 1521 -64 1897
rect 0 1521 34 1897
rect 98 1521 132 1897
rect 196 1521 230 1897
rect 294 1521 328 1897
rect 622 2157 656 2533
rect 720 2157 754 2533
rect 818 2157 852 2533
rect 916 2157 950 2533
rect 1014 2157 1048 2533
rect 1112 2157 1146 2533
rect 1210 2157 1244 2533
rect 1308 2157 1342 2533
rect 1406 2157 1440 2533
rect 1504 2157 1538 2533
rect 1602 2157 1636 2533
rect 1700 2157 1734 2533
rect 1798 2157 1832 2533
rect 1896 2157 1930 2533
rect 1994 2157 2028 2533
rect 2092 2157 2126 2533
rect 622 1521 656 1897
rect 720 1521 754 1897
rect 818 1521 852 1897
rect 916 1521 950 1897
rect 1014 1521 1048 1897
rect 1112 1521 1146 1897
rect 1210 1521 1244 1897
rect 1308 1521 1342 1897
rect 1406 1521 1440 1897
rect 1504 1521 1538 1897
rect 1602 1521 1636 1897
rect 1700 1521 1734 1897
rect 1798 1521 1832 1897
rect 1896 1521 1930 1897
rect 1994 1521 2028 1897
rect 2092 1521 2126 1897
rect 2424 1505 2458 1881
rect 2582 1505 2616 1881
rect 2740 1505 2774 1881
rect 2898 1505 2932 1881
rect 3056 1505 3090 1881
rect 3214 1505 3248 1881
rect 3372 1505 3406 1881
rect 3530 1505 3564 1881
rect 3688 1505 3722 1881
rect 3846 1505 3880 1881
rect 4004 1505 4038 1881
rect -1176 -4913 -1142 -4537
rect -1078 -4913 -1044 -4537
rect -980 -4913 -946 -4537
rect -882 -4913 -848 -4537
rect -784 -4913 -750 -4537
rect -686 -4913 -652 -4537
rect -588 -4913 -554 -4537
rect -490 -4913 -456 -4537
rect -392 -4913 -358 -4537
rect -294 -4913 -260 -4537
rect -196 -4913 -162 -4537
rect -98 -4913 -64 -4537
rect 0 -4913 34 -4537
rect 98 -4913 132 -4537
rect 196 -4913 230 -4537
rect 294 -4913 328 -4537
rect -1176 -5549 -1142 -5173
rect -1078 -5549 -1044 -5173
rect -980 -5549 -946 -5173
rect -882 -5549 -848 -5173
rect -784 -5549 -750 -5173
rect -686 -5549 -652 -5173
rect -588 -5549 -554 -5173
rect -490 -5549 -456 -5173
rect -392 -5549 -358 -5173
rect -294 -5549 -260 -5173
rect -196 -5549 -162 -5173
rect -98 -5549 -64 -5173
rect 0 -5549 34 -5173
rect 98 -5549 132 -5173
rect 196 -5549 230 -5173
rect 294 -5549 328 -5173
rect 622 -4913 656 -4537
rect 720 -4913 754 -4537
rect 818 -4913 852 -4537
rect 916 -4913 950 -4537
rect 1014 -4913 1048 -4537
rect 1112 -4913 1146 -4537
rect 1210 -4913 1244 -4537
rect 1308 -4913 1342 -4537
rect 1406 -4913 1440 -4537
rect 1504 -4913 1538 -4537
rect 1602 -4913 1636 -4537
rect 1700 -4913 1734 -4537
rect 1798 -4913 1832 -4537
rect 1896 -4913 1930 -4537
rect 1994 -4913 2028 -4537
rect 2092 -4913 2126 -4537
rect 622 -5549 656 -5173
rect 720 -5549 754 -5173
rect 818 -5549 852 -5173
rect 916 -5549 950 -5173
rect 1014 -5549 1048 -5173
rect 1112 -5549 1146 -5173
rect 1210 -5549 1244 -5173
rect 1308 -5549 1342 -5173
rect 1406 -5549 1440 -5173
rect 1504 -5549 1538 -5173
rect 1602 -5549 1636 -5173
rect 1700 -5549 1734 -5173
rect 1798 -5549 1832 -5173
rect 1896 -5549 1930 -5173
rect 1994 -5549 2028 -5173
rect 2092 -5549 2126 -5173
rect 2424 -5565 2458 -5189
rect 2582 -5565 2616 -5189
rect 2740 -5565 2774 -5189
rect 2898 -5565 2932 -5189
rect 3056 -5565 3090 -5189
rect 3214 -5565 3248 -5189
rect 3372 -5565 3406 -5189
rect 3530 -5565 3564 -5189
rect 3688 -5565 3722 -5189
rect 3846 -5565 3880 -5189
rect 4004 -5565 4038 -5189
rect 6330 -10299 6364 -10223
rect 6588 -10299 6622 -10223
<< psubdiff >>
rect -1290 1218 -1194 1252
rect 1326 1218 1422 1252
rect -1290 1156 -1256 1218
rect 1388 1156 1422 1218
rect -1290 -80 -1256 -18
rect 1388 -80 1422 -18
rect -1290 -114 -1194 -80
rect 1326 -114 1422 -80
rect -1290 -226 -1194 -192
rect 1326 -226 1422 -192
rect -1290 -288 -1256 -226
rect 1388 -288 1422 -226
rect -1290 -1524 -1256 -1462
rect 2370 898 2466 932
rect 4006 898 4102 932
rect 2370 836 2404 898
rect 4068 836 4102 898
rect 2370 -400 2404 -338
rect 4068 -400 4102 -338
rect 2370 -434 2466 -400
rect 4006 -434 4102 -400
rect 1388 -1524 1422 -1462
rect -1290 -1558 -1194 -1524
rect 1326 -1558 1422 -1524
rect 1500 -880 1596 -846
rect 2818 -880 2914 -846
rect 1500 -942 1534 -880
rect 2880 -942 2914 -880
rect 1500 -1560 1534 -1498
rect 2880 -1560 2914 -1498
rect 1500 -1594 1596 -1560
rect 2818 -1594 2914 -1560
rect -1310 -1646 -1214 -1612
rect 1256 -1646 1352 -1612
rect -1310 -1708 -1276 -1646
rect 1318 -1708 1352 -1646
rect -1310 -4180 -1276 -4118
rect 1500 -1700 1596 -1666
rect 3214 -1700 3310 -1666
rect 1500 -1762 1534 -1700
rect 3276 -1762 3310 -1700
rect 1500 -2380 1534 -2318
rect 3276 -2380 3310 -2318
rect 1500 -2414 1596 -2380
rect 3214 -2414 3310 -2380
rect 1318 -4180 1352 -4118
rect -1310 -4214 -1214 -4180
rect 1256 -4214 1352 -4180
rect -1290 -5852 -1194 -5818
rect 1326 -5852 1422 -5818
rect -1290 -5914 -1256 -5852
rect 1388 -5914 1422 -5852
rect -1290 -7150 -1256 -7088
rect 1388 -7150 1422 -7088
rect -1290 -7184 -1194 -7150
rect 1326 -7184 1422 -7150
rect -1290 -7296 -1194 -7262
rect 1326 -7296 1422 -7262
rect -1290 -7358 -1256 -7296
rect 1388 -7358 1422 -7296
rect -1290 -8594 -1256 -8532
rect 2370 -6172 2466 -6138
rect 4006 -6172 4102 -6138
rect 2370 -6234 2404 -6172
rect 4068 -6234 4102 -6172
rect 2370 -7470 2404 -7408
rect 4068 -7470 4102 -7408
rect 2370 -7504 2466 -7470
rect 4006 -7504 4102 -7470
rect 1388 -8594 1422 -8532
rect -1290 -8628 -1194 -8594
rect 1326 -8628 1422 -8594
rect 1500 -7950 1596 -7916
rect 2818 -7950 2914 -7916
rect 1500 -8012 1534 -7950
rect 2880 -8012 2914 -7950
rect 1500 -8630 1534 -8568
rect 2880 -8630 2914 -8568
rect 1500 -8664 1596 -8630
rect 2818 -8664 2914 -8630
rect 3396 -7950 3492 -7916
rect 4714 -7950 4810 -7916
rect 3396 -8012 3430 -7950
rect 4776 -8012 4810 -7950
rect 3396 -8630 3430 -8568
rect 4776 -8630 4810 -8568
rect 3396 -8664 3492 -8630
rect 4714 -8664 4810 -8630
rect -1310 -8716 -1214 -8682
rect 1256 -8716 1352 -8682
rect -1310 -8778 -1276 -8716
rect 1318 -8778 1352 -8716
rect -1310 -11250 -1276 -11188
rect 1500 -8770 1596 -8736
rect 3214 -8770 3310 -8736
rect 1500 -8832 1534 -8770
rect 3276 -8832 3310 -8770
rect 1500 -9450 1534 -9388
rect 3276 -9450 3310 -9388
rect 1500 -9484 1596 -9450
rect 3214 -9484 3310 -9450
rect 3396 -8770 3492 -8736
rect 5110 -8770 5206 -8736
rect 3396 -8832 3430 -8770
rect 5172 -8832 5206 -8770
rect 3396 -9450 3430 -9388
rect 5172 -9450 5206 -9388
rect 3396 -9484 3492 -9450
rect 5110 -9484 5206 -9450
rect 5346 -8770 5442 -8736
rect 5992 -8770 6088 -8736
rect 5346 -8832 5380 -8770
rect 6054 -8832 6088 -8770
rect 5346 -9450 5380 -9388
rect 6054 -9450 6088 -9388
rect 5346 -9484 5442 -9450
rect 5992 -9484 6088 -9450
rect 1486 -9764 1582 -9730
rect 5884 -9764 5980 -9730
rect 1486 -9853 1520 -9764
rect 5946 -9853 5980 -9764
rect 1486 -11080 1520 -10991
rect 5946 -11080 5980 -10991
rect 6216 -10630 6312 -10596
rect 6640 -10630 6736 -10596
rect 6216 -10692 6250 -10630
rect 6702 -10692 6736 -10630
rect 6216 -11010 6250 -10948
rect 6702 -11010 6736 -10948
rect 6216 -11044 6312 -11010
rect 6640 -11044 6736 -11010
rect 1486 -11114 1609 -11080
rect 5857 -11114 5980 -11080
rect 1318 -11250 1352 -11188
rect -1310 -11284 -1214 -11250
rect 1256 -11284 1352 -11250
<< nsubdiff >>
rect -1290 2694 -1194 2728
rect 346 2694 442 2728
rect -1290 2632 -1256 2694
rect 408 2632 442 2694
rect -1290 1360 -1256 1422
rect 408 1360 442 1422
rect -1290 1326 -1194 1360
rect 346 1326 442 1360
rect 508 2694 604 2728
rect 2144 2694 2240 2728
rect 508 2632 542 2694
rect 2206 2632 2240 2694
rect 508 1360 542 1422
rect 2206 1360 2240 1422
rect 508 1326 604 1360
rect 2144 1326 2240 1360
rect 2310 2042 2406 2076
rect 4056 2042 4152 2076
rect 2310 1980 2344 2042
rect 4118 1980 4152 2042
rect 2310 1344 2344 1406
rect 4118 1344 4152 1406
rect 2310 1310 2406 1344
rect 4056 1310 4152 1344
rect 2051 1233 4417 1253
rect 2051 1199 2131 1233
rect 4337 1199 4417 1233
rect 2051 1179 4417 1199
rect 2051 1173 2125 1179
rect 2051 -673 2071 1173
rect 2105 -673 2125 1173
rect 4343 1173 4417 1179
rect 2051 -679 2125 -673
rect 4343 -673 4363 1173
rect 4397 -673 4417 1173
rect 4343 -679 4417 -673
rect 2051 -699 4417 -679
rect 2051 -733 2131 -699
rect 4337 -733 4417 -699
rect 2051 -753 4417 -733
rect -1290 -4376 -1194 -4342
rect 346 -4376 442 -4342
rect -1290 -4438 -1256 -4376
rect 408 -4438 442 -4376
rect -1290 -5710 -1256 -5648
rect 408 -5710 442 -5648
rect -1290 -5744 -1194 -5710
rect 346 -5744 442 -5710
rect 508 -4376 604 -4342
rect 2144 -4376 2240 -4342
rect 508 -4438 542 -4376
rect 2206 -4438 2240 -4376
rect 508 -5710 542 -5648
rect 2206 -5710 2240 -5648
rect 508 -5744 604 -5710
rect 2144 -5744 2240 -5710
rect 2310 -5028 2406 -4994
rect 4056 -5028 4152 -4994
rect 2310 -5090 2344 -5028
rect 4118 -5090 4152 -5028
rect 2310 -5726 2344 -5664
rect 4118 -5726 4152 -5664
rect 2310 -5760 2406 -5726
rect 4056 -5760 4152 -5726
rect 2051 -5837 4417 -5817
rect 2051 -5871 2131 -5837
rect 4337 -5871 4417 -5837
rect 2051 -5891 4417 -5871
rect 2051 -5897 2125 -5891
rect 2051 -7743 2071 -5897
rect 2105 -7743 2125 -5897
rect 4343 -5897 4417 -5891
rect 2051 -7749 2125 -7743
rect 4343 -7743 4363 -5897
rect 4397 -7743 4417 -5897
rect 4343 -7749 4417 -7743
rect 2051 -7769 4417 -7749
rect 2051 -7803 2131 -7769
rect 4337 -7803 4417 -7769
rect 2051 -7823 4417 -7803
rect 1596 -9946 1693 -9922
rect 1596 -10898 1608 -9946
rect 1642 -10898 1693 -9946
rect 1596 -10922 1693 -10898
rect 2093 -9946 2190 -9922
rect 2093 -10898 2144 -9946
rect 2178 -10898 2190 -9946
rect 2093 -10922 2190 -10898
rect 2516 -9946 2613 -9922
rect 2516 -10898 2528 -9946
rect 2562 -10898 2613 -9946
rect 2516 -10922 2613 -10898
rect 3013 -9946 3110 -9922
rect 3013 -10898 3064 -9946
rect 3098 -10898 3110 -9946
rect 3013 -10922 3110 -10898
rect 3436 -9946 3533 -9922
rect 3436 -10898 3448 -9946
rect 3482 -10898 3533 -9946
rect 3436 -10922 3533 -10898
rect 3933 -9946 4030 -9922
rect 3933 -10898 3984 -9946
rect 4018 -10898 4030 -9946
rect 3933 -10922 4030 -10898
rect 4356 -9946 4453 -9922
rect 4356 -10898 4368 -9946
rect 4402 -10898 4453 -9946
rect 4356 -10922 4453 -10898
rect 4853 -9946 4950 -9922
rect 4853 -10898 4904 -9946
rect 4938 -10898 4950 -9946
rect 4853 -10922 4950 -10898
rect 5276 -9946 5373 -9922
rect 5276 -10898 5288 -9946
rect 5322 -10898 5373 -9946
rect 5276 -10922 5373 -10898
rect 5773 -9946 5870 -9922
rect 5773 -10898 5824 -9946
rect 5858 -10898 5870 -9946
rect 5773 -10922 5870 -10898
rect 6216 -10062 6312 -10028
rect 6640 -10062 6736 -10028
rect 6216 -10124 6250 -10062
rect 6702 -10124 6736 -10062
rect 6216 -10460 6250 -10398
rect 6702 -10460 6736 -10398
rect 6216 -10494 6312 -10460
rect 6640 -10494 6736 -10460
<< psubdiffcont >>
rect -1194 1218 1326 1252
rect -1290 -18 -1256 1156
rect 1388 -18 1422 1156
rect -1194 -114 1326 -80
rect -1194 -226 1326 -192
rect -1290 -1462 -1256 -288
rect 1388 -1462 1422 -288
rect 2466 898 4006 932
rect 2370 -338 2404 836
rect 4068 -338 4102 836
rect 2466 -434 4006 -400
rect -1194 -1558 1326 -1524
rect 1596 -880 2818 -846
rect 1500 -1498 1534 -942
rect 2880 -1498 2914 -942
rect 1596 -1594 2818 -1560
rect -1214 -1646 1256 -1612
rect -1310 -4118 -1276 -1708
rect 1318 -4118 1352 -1708
rect 1596 -1700 3214 -1666
rect 1500 -2318 1534 -1762
rect 3276 -2318 3310 -1762
rect 1596 -2414 3214 -2380
rect -1214 -4214 1256 -4180
rect -1194 -5852 1326 -5818
rect -1290 -7088 -1256 -5914
rect 1388 -7088 1422 -5914
rect -1194 -7184 1326 -7150
rect -1194 -7296 1326 -7262
rect -1290 -8532 -1256 -7358
rect 1388 -8532 1422 -7358
rect 2466 -6172 4006 -6138
rect 2370 -7408 2404 -6234
rect 4068 -7408 4102 -6234
rect 2466 -7504 4006 -7470
rect -1194 -8628 1326 -8594
rect 1596 -7950 2818 -7916
rect 1500 -8568 1534 -8012
rect 2880 -8568 2914 -8012
rect 1596 -8664 2818 -8630
rect 3492 -7950 4714 -7916
rect 3396 -8568 3430 -8012
rect 4776 -8568 4810 -8012
rect 3492 -8664 4714 -8630
rect -1214 -8716 1256 -8682
rect -1310 -11188 -1276 -8778
rect 1318 -11188 1352 -8778
rect 1596 -8770 3214 -8736
rect 1500 -9388 1534 -8832
rect 3276 -9388 3310 -8832
rect 1596 -9484 3214 -9450
rect 3492 -8770 5110 -8736
rect 3396 -9388 3430 -8832
rect 5172 -9388 5206 -8832
rect 3492 -9484 5110 -9450
rect 5442 -8770 5992 -8736
rect 5346 -9388 5380 -8832
rect 6054 -9388 6088 -8832
rect 5442 -9484 5992 -9450
rect 1582 -9764 5884 -9730
rect 1486 -10991 1520 -9853
rect 5946 -10991 5980 -9853
rect 6312 -10630 6640 -10596
rect 6216 -10948 6250 -10692
rect 6702 -10948 6736 -10692
rect 6312 -11044 6640 -11010
rect 1609 -11114 5857 -11080
rect -1214 -11284 1256 -11250
<< nsubdiffcont >>
rect -1194 2694 346 2728
rect -1290 1422 -1256 2632
rect 408 1422 442 2632
rect -1194 1326 346 1360
rect 604 2694 2144 2728
rect 508 1422 542 2632
rect 2206 1422 2240 2632
rect 604 1326 2144 1360
rect 2406 2042 4056 2076
rect 2310 1406 2344 1980
rect 4118 1406 4152 1980
rect 2406 1310 4056 1344
rect 2131 1199 4337 1233
rect 2071 -673 2105 1173
rect 4363 -673 4397 1173
rect 2131 -733 4337 -699
rect -1194 -4376 346 -4342
rect -1290 -5648 -1256 -4438
rect 408 -5648 442 -4438
rect -1194 -5744 346 -5710
rect 604 -4376 2144 -4342
rect 508 -5648 542 -4438
rect 2206 -5648 2240 -4438
rect 604 -5744 2144 -5710
rect 2406 -5028 4056 -4994
rect 2310 -5664 2344 -5090
rect 4118 -5664 4152 -5090
rect 2406 -5760 4056 -5726
rect 2131 -5871 4337 -5837
rect 2071 -7743 2105 -5897
rect 4363 -7743 4397 -5897
rect 2131 -7803 4337 -7769
rect 1608 -10898 1642 -9946
rect 2144 -10898 2178 -9946
rect 2528 -10898 2562 -9946
rect 3064 -10898 3098 -9946
rect 3448 -10898 3482 -9946
rect 3984 -10898 4018 -9946
rect 4368 -10898 4402 -9946
rect 4904 -10898 4938 -9946
rect 5288 -10898 5322 -9946
rect 5824 -10898 5858 -9946
rect 6312 -10062 6640 -10028
rect 6216 -10398 6250 -10124
rect 6702 -10398 6736 -10124
rect 6312 -10494 6640 -10460
<< poly >>
rect -1143 2626 295 2642
rect -1143 2592 -1127 2626
rect -1093 2592 -1029 2626
rect -995 2592 -931 2626
rect -897 2592 -833 2626
rect -799 2592 -735 2626
rect -701 2592 -637 2626
rect -603 2592 -539 2626
rect -505 2592 -441 2626
rect -407 2592 -343 2626
rect -309 2592 -245 2626
rect -211 2592 -147 2626
rect -113 2592 -49 2626
rect -15 2592 49 2626
rect 83 2592 147 2626
rect 181 2592 245 2626
rect 279 2592 295 2626
rect -1143 2576 295 2592
rect -1130 2545 -1090 2576
rect -1032 2545 -992 2576
rect -934 2545 -894 2576
rect -836 2545 -796 2576
rect -738 2545 -698 2576
rect -640 2545 -600 2576
rect -542 2545 -502 2576
rect -444 2545 -404 2576
rect -346 2545 -306 2576
rect -248 2545 -208 2576
rect -150 2545 -110 2576
rect -52 2545 -12 2576
rect 46 2545 86 2576
rect 144 2545 184 2576
rect 242 2545 282 2576
rect -1130 2114 -1090 2145
rect -1032 2114 -992 2145
rect -934 2114 -894 2145
rect -836 2114 -796 2145
rect -738 2114 -698 2145
rect -640 2114 -600 2145
rect -542 2114 -502 2145
rect -444 2114 -404 2145
rect -346 2114 -306 2145
rect -248 2114 -208 2145
rect -150 2114 -110 2145
rect -52 2114 -12 2145
rect 46 2114 86 2145
rect 144 2114 184 2145
rect 242 2114 282 2145
rect -1143 2098 295 2114
rect -1143 2064 -1127 2098
rect -1093 2064 -1029 2098
rect -995 2064 -931 2098
rect -897 2064 -833 2098
rect -799 2064 -735 2098
rect -701 2064 -637 2098
rect -603 2064 -539 2098
rect -505 2064 -441 2098
rect -407 2064 -343 2098
rect -309 2064 -245 2098
rect -211 2064 -147 2098
rect -113 2064 -49 2098
rect -15 2064 49 2098
rect 83 2064 147 2098
rect 181 2064 245 2098
rect 279 2064 295 2098
rect -1143 2048 295 2064
rect -1143 1990 295 2006
rect -1143 1956 -1127 1990
rect -1093 1956 -1029 1990
rect -995 1956 -931 1990
rect -897 1956 -833 1990
rect -799 1956 -735 1990
rect -701 1956 -637 1990
rect -603 1956 -539 1990
rect -505 1956 -441 1990
rect -407 1956 -343 1990
rect -309 1956 -245 1990
rect -211 1956 -147 1990
rect -113 1956 -49 1990
rect -15 1956 49 1990
rect 83 1956 147 1990
rect 181 1956 245 1990
rect 279 1956 295 1990
rect -1143 1940 295 1956
rect -1130 1909 -1090 1940
rect -1032 1909 -992 1940
rect -934 1909 -894 1940
rect -836 1909 -796 1940
rect -738 1909 -698 1940
rect -640 1909 -600 1940
rect -542 1909 -502 1940
rect -444 1909 -404 1940
rect -346 1909 -306 1940
rect -248 1909 -208 1940
rect -150 1909 -110 1940
rect -52 1909 -12 1940
rect 46 1909 86 1940
rect 144 1909 184 1940
rect 242 1909 282 1940
rect -1130 1478 -1090 1509
rect -1032 1478 -992 1509
rect -934 1478 -894 1509
rect -836 1478 -796 1509
rect -738 1478 -698 1509
rect -640 1478 -600 1509
rect -542 1478 -502 1509
rect -444 1478 -404 1509
rect -346 1478 -306 1509
rect -248 1478 -208 1509
rect -150 1478 -110 1509
rect -52 1478 -12 1509
rect 46 1478 86 1509
rect 144 1478 184 1509
rect 242 1478 282 1509
rect -1143 1462 295 1478
rect -1143 1428 -1127 1462
rect -1093 1428 -1029 1462
rect -995 1428 -931 1462
rect -897 1428 -833 1462
rect -799 1428 -735 1462
rect -701 1428 -637 1462
rect -603 1428 -539 1462
rect -505 1428 -441 1462
rect -407 1428 -343 1462
rect -309 1428 -245 1462
rect -211 1428 -147 1462
rect -113 1428 -49 1462
rect -15 1428 49 1462
rect 83 1428 147 1462
rect 181 1428 245 1462
rect 279 1428 295 1462
rect -1143 1412 295 1428
rect 655 2626 2093 2642
rect 655 2592 671 2626
rect 705 2592 769 2626
rect 803 2592 867 2626
rect 901 2592 965 2626
rect 999 2592 1063 2626
rect 1097 2592 1161 2626
rect 1195 2592 1259 2626
rect 1293 2592 1357 2626
rect 1391 2592 1455 2626
rect 1489 2592 1553 2626
rect 1587 2592 1651 2626
rect 1685 2592 1749 2626
rect 1783 2592 1847 2626
rect 1881 2592 1945 2626
rect 1979 2592 2043 2626
rect 2077 2592 2093 2626
rect 655 2576 2093 2592
rect 668 2545 708 2576
rect 766 2545 806 2576
rect 864 2545 904 2576
rect 962 2545 1002 2576
rect 1060 2545 1100 2576
rect 1158 2545 1198 2576
rect 1256 2545 1296 2576
rect 1354 2545 1394 2576
rect 1452 2545 1492 2576
rect 1550 2545 1590 2576
rect 1648 2545 1688 2576
rect 1746 2545 1786 2576
rect 1844 2545 1884 2576
rect 1942 2545 1982 2576
rect 2040 2545 2080 2576
rect 668 2114 708 2145
rect 766 2114 806 2145
rect 864 2114 904 2145
rect 962 2114 1002 2145
rect 1060 2114 1100 2145
rect 1158 2114 1198 2145
rect 1256 2114 1296 2145
rect 1354 2114 1394 2145
rect 1452 2114 1492 2145
rect 1550 2114 1590 2145
rect 1648 2114 1688 2145
rect 1746 2114 1786 2145
rect 1844 2114 1884 2145
rect 1942 2114 1982 2145
rect 2040 2114 2080 2145
rect 655 2098 2093 2114
rect 655 2064 671 2098
rect 705 2064 769 2098
rect 803 2064 867 2098
rect 901 2064 965 2098
rect 999 2064 1063 2098
rect 1097 2064 1161 2098
rect 1195 2064 1259 2098
rect 1293 2064 1357 2098
rect 1391 2064 1455 2098
rect 1489 2064 1553 2098
rect 1587 2064 1651 2098
rect 1685 2064 1749 2098
rect 1783 2064 1847 2098
rect 1881 2064 1945 2098
rect 1979 2064 2043 2098
rect 2077 2064 2093 2098
rect 655 2048 2093 2064
rect 655 1990 2093 2006
rect 655 1956 671 1990
rect 705 1956 769 1990
rect 803 1956 867 1990
rect 901 1956 965 1990
rect 999 1956 1063 1990
rect 1097 1956 1161 1990
rect 1195 1956 1259 1990
rect 1293 1956 1357 1990
rect 1391 1956 1455 1990
rect 1489 1956 1553 1990
rect 1587 1956 1651 1990
rect 1685 1956 1749 1990
rect 1783 1956 1847 1990
rect 1881 1956 1945 1990
rect 1979 1956 2043 1990
rect 2077 1956 2093 1990
rect 655 1940 2093 1956
rect 668 1909 708 1940
rect 766 1909 806 1940
rect 864 1909 904 1940
rect 962 1909 1002 1940
rect 1060 1909 1100 1940
rect 1158 1909 1198 1940
rect 1256 1909 1296 1940
rect 1354 1909 1394 1940
rect 1452 1909 1492 1940
rect 1550 1909 1590 1940
rect 1648 1909 1688 1940
rect 1746 1909 1786 1940
rect 1844 1909 1884 1940
rect 1942 1909 1982 1940
rect 2040 1909 2080 1940
rect 668 1478 708 1509
rect 766 1478 806 1509
rect 864 1478 904 1509
rect 962 1478 1002 1509
rect 1060 1478 1100 1509
rect 1158 1478 1198 1509
rect 1256 1478 1296 1509
rect 1354 1478 1394 1509
rect 1452 1478 1492 1509
rect 1550 1478 1590 1509
rect 1648 1478 1688 1509
rect 1746 1478 1786 1509
rect 1844 1478 1884 1509
rect 1942 1478 1982 1509
rect 2040 1478 2080 1509
rect 655 1462 2093 1478
rect 655 1428 671 1462
rect 705 1428 769 1462
rect 803 1428 867 1462
rect 901 1428 965 1462
rect 999 1428 1063 1462
rect 1097 1428 1161 1462
rect 1195 1428 1259 1462
rect 1293 1428 1357 1462
rect 1391 1428 1455 1462
rect 1489 1428 1553 1462
rect 1587 1428 1651 1462
rect 1685 1428 1749 1462
rect 1783 1428 1847 1462
rect 1881 1428 1945 1462
rect 1979 1428 2043 1462
rect 2077 1428 2093 1462
rect 655 1412 2093 1428
rect 2470 1974 2570 1990
rect 2470 1940 2486 1974
rect 2554 1940 2570 1974
rect 2470 1893 2570 1940
rect 2628 1974 2728 1990
rect 2628 1940 2644 1974
rect 2712 1940 2728 1974
rect 2628 1893 2728 1940
rect 2786 1974 2886 1990
rect 2786 1940 2802 1974
rect 2870 1940 2886 1974
rect 2786 1893 2886 1940
rect 2944 1974 3044 1990
rect 2944 1940 2960 1974
rect 3028 1940 3044 1974
rect 2944 1893 3044 1940
rect 3102 1974 3202 1990
rect 3102 1940 3118 1974
rect 3186 1940 3202 1974
rect 3102 1893 3202 1940
rect 3260 1974 3360 1990
rect 3260 1940 3276 1974
rect 3344 1940 3360 1974
rect 3260 1893 3360 1940
rect 3418 1974 3518 1990
rect 3418 1940 3434 1974
rect 3502 1940 3518 1974
rect 3418 1893 3518 1940
rect 3576 1974 3676 1990
rect 3576 1940 3592 1974
rect 3660 1940 3676 1974
rect 3576 1893 3676 1940
rect 3734 1974 3834 1990
rect 3734 1940 3750 1974
rect 3818 1940 3834 1974
rect 3734 1893 3834 1940
rect 3892 1974 3992 1990
rect 3892 1940 3908 1974
rect 3976 1940 3992 1974
rect 3892 1893 3992 1940
rect 2470 1446 2570 1493
rect 2470 1412 2486 1446
rect 2554 1412 2570 1446
rect 2470 1396 2570 1412
rect 2628 1446 2728 1493
rect 2628 1412 2644 1446
rect 2712 1412 2728 1446
rect 2628 1396 2728 1412
rect 2786 1446 2886 1493
rect 2786 1412 2802 1446
rect 2870 1412 2886 1446
rect 2786 1396 2886 1412
rect 2944 1446 3044 1493
rect 2944 1412 2960 1446
rect 3028 1412 3044 1446
rect 2944 1396 3044 1412
rect 3102 1446 3202 1493
rect 3102 1412 3118 1446
rect 3186 1412 3202 1446
rect 3102 1396 3202 1412
rect 3260 1446 3360 1493
rect 3260 1412 3276 1446
rect 3344 1412 3360 1446
rect 3260 1396 3360 1412
rect 3418 1446 3518 1493
rect 3418 1412 3434 1446
rect 3502 1412 3518 1446
rect 3418 1396 3518 1412
rect 3576 1446 3676 1493
rect 3576 1412 3592 1446
rect 3660 1412 3676 1446
rect 3576 1396 3676 1412
rect 3734 1446 3834 1493
rect 3734 1412 3750 1446
rect 3818 1412 3834 1446
rect 3734 1396 3834 1412
rect 3892 1446 3992 1493
rect 3892 1412 3908 1446
rect 3976 1412 3992 1446
rect 3892 1396 3992 1412
rect -1144 1150 1275 1166
rect -1144 1116 -1127 1150
rect -1093 1116 -1030 1150
rect -996 1116 -931 1150
rect -897 1116 -834 1150
rect -800 1116 -735 1150
rect -701 1116 -638 1150
rect -604 1116 -539 1150
rect -505 1116 -442 1150
rect -408 1116 -343 1150
rect -309 1116 -246 1150
rect -212 1116 -147 1150
rect -113 1116 -50 1150
rect -16 1116 49 1150
rect 83 1116 146 1150
rect 180 1116 245 1150
rect 279 1116 342 1150
rect 376 1116 441 1150
rect 475 1116 538 1150
rect 572 1116 637 1150
rect 671 1116 734 1150
rect 768 1116 833 1150
rect 867 1116 930 1150
rect 964 1116 1029 1150
rect 1063 1116 1126 1150
rect 1160 1116 1225 1150
rect 1259 1116 1275 1150
rect -1144 1100 1275 1116
rect -1130 1078 -1090 1100
rect -1032 1078 -992 1100
rect -934 1078 -894 1100
rect -836 1078 -796 1100
rect -738 1078 -698 1100
rect -640 1078 -600 1100
rect -542 1078 -502 1100
rect -444 1078 -404 1100
rect -346 1078 -306 1100
rect -248 1078 -208 1100
rect -150 1078 -110 1100
rect -52 1078 -12 1100
rect 46 1078 86 1100
rect 144 1078 184 1100
rect 242 1078 282 1100
rect 340 1078 380 1100
rect 438 1078 478 1100
rect 536 1078 576 1100
rect 634 1078 674 1100
rect 732 1078 772 1100
rect 830 1078 870 1100
rect 928 1078 968 1100
rect 1026 1078 1066 1100
rect 1124 1078 1164 1100
rect 1222 1078 1262 1100
rect -1130 656 -1090 678
rect -1032 656 -992 678
rect -934 656 -894 678
rect -836 656 -796 678
rect -738 656 -698 678
rect -640 656 -600 678
rect -542 656 -502 678
rect -444 656 -404 678
rect -346 656 -306 678
rect -248 656 -208 678
rect -150 656 -110 678
rect -52 656 -12 678
rect 46 656 86 678
rect 144 656 184 678
rect 242 656 282 678
rect 340 656 380 678
rect 438 656 478 678
rect 536 656 576 678
rect 634 656 674 678
rect 732 656 772 678
rect 830 656 870 678
rect 928 656 968 678
rect 1026 656 1066 678
rect 1124 656 1164 678
rect 1222 656 1262 678
rect -1144 640 1274 656
rect -1144 606 -1128 640
rect -1094 606 -1029 640
rect -995 606 -932 640
rect -898 606 -833 640
rect -799 606 -736 640
rect -702 606 -637 640
rect -603 606 -540 640
rect -506 606 -441 640
rect -407 606 -344 640
rect -310 606 -245 640
rect -211 606 -148 640
rect -114 606 -49 640
rect -15 606 48 640
rect 82 606 147 640
rect 181 606 244 640
rect 278 606 343 640
rect 377 606 440 640
rect 474 606 539 640
rect 573 606 636 640
rect 670 606 735 640
rect 769 606 832 640
rect 866 606 931 640
rect 965 606 1028 640
rect 1062 606 1127 640
rect 1161 606 1224 640
rect 1258 606 1274 640
rect -1144 590 1274 606
rect -1143 532 1275 548
rect -1143 498 -1127 532
rect -1093 498 -1029 532
rect -995 498 -931 532
rect -897 498 -833 532
rect -799 498 -735 532
rect -701 498 -637 532
rect -603 498 -539 532
rect -505 498 -441 532
rect -407 498 -343 532
rect -309 498 -245 532
rect -211 498 -147 532
rect -113 498 -49 532
rect -15 498 49 532
rect 83 498 147 532
rect 181 498 245 532
rect 279 498 343 532
rect 377 498 441 532
rect 475 498 539 532
rect 573 498 637 532
rect 671 498 735 532
rect 769 498 833 532
rect 867 498 931 532
rect 965 498 1029 532
rect 1063 498 1127 532
rect 1161 498 1225 532
rect 1259 498 1275 532
rect -1143 482 1275 498
rect -1130 460 -1090 482
rect -1032 460 -992 482
rect -934 460 -894 482
rect -836 460 -796 482
rect -738 460 -698 482
rect -640 460 -600 482
rect -542 460 -502 482
rect -444 460 -404 482
rect -346 460 -306 482
rect -248 460 -208 482
rect -150 460 -110 482
rect -52 460 -12 482
rect 46 460 86 482
rect 144 460 184 482
rect 242 460 282 482
rect 340 460 380 482
rect 438 460 478 482
rect 536 460 576 482
rect 634 460 674 482
rect 732 460 772 482
rect 830 460 870 482
rect 928 460 968 482
rect 1026 460 1066 482
rect 1124 460 1164 482
rect 1222 460 1262 482
rect -1130 38 -1090 60
rect -1032 38 -992 60
rect -934 38 -894 60
rect -836 38 -796 60
rect -738 38 -698 60
rect -640 38 -600 60
rect -542 38 -502 60
rect -444 38 -404 60
rect -346 38 -306 60
rect -248 38 -208 60
rect -150 38 -110 60
rect -52 38 -12 60
rect 46 38 86 60
rect 144 38 184 60
rect 242 38 282 60
rect 340 38 380 60
rect 438 38 478 60
rect 536 38 576 60
rect 634 38 674 60
rect 732 38 772 60
rect 830 38 870 60
rect 928 38 968 60
rect 1026 38 1066 60
rect 1124 38 1164 60
rect 1222 38 1262 60
rect -1143 22 1275 38
rect -1143 -12 -1127 22
rect -1093 -12 -1029 22
rect -995 -12 -931 22
rect -897 -12 -833 22
rect -799 -12 -735 22
rect -701 -12 -637 22
rect -603 -12 -539 22
rect -505 -12 -441 22
rect -407 -12 -343 22
rect -309 -12 -245 22
rect -211 -12 -147 22
rect -113 -12 -49 22
rect -15 -12 49 22
rect 83 -12 147 22
rect 181 -12 245 22
rect 279 -12 343 22
rect 377 -12 441 22
rect 475 -12 539 22
rect 573 -12 637 22
rect 671 -12 735 22
rect 769 -12 833 22
rect 867 -12 931 22
rect 965 -12 1029 22
rect 1063 -12 1127 22
rect 1161 -12 1225 22
rect 1259 -12 1275 22
rect -1143 -28 1275 -12
rect -1144 -294 1275 -278
rect -1144 -328 -1127 -294
rect -1093 -328 -1030 -294
rect -996 -328 -931 -294
rect -897 -328 -834 -294
rect -800 -328 -735 -294
rect -701 -328 -638 -294
rect -604 -328 -539 -294
rect -505 -328 -442 -294
rect -408 -328 -343 -294
rect -309 -328 -246 -294
rect -212 -328 -147 -294
rect -113 -328 -50 -294
rect -16 -328 49 -294
rect 83 -328 146 -294
rect 180 -328 245 -294
rect 279 -328 342 -294
rect 376 -328 441 -294
rect 475 -328 538 -294
rect 572 -328 637 -294
rect 671 -328 734 -294
rect 768 -328 833 -294
rect 867 -328 930 -294
rect 964 -328 1029 -294
rect 1063 -328 1126 -294
rect 1160 -328 1225 -294
rect 1259 -328 1275 -294
rect -1144 -344 1275 -328
rect -1130 -366 -1090 -344
rect -1032 -366 -992 -344
rect -934 -366 -894 -344
rect -836 -366 -796 -344
rect -738 -366 -698 -344
rect -640 -366 -600 -344
rect -542 -366 -502 -344
rect -444 -366 -404 -344
rect -346 -366 -306 -344
rect -248 -366 -208 -344
rect -150 -366 -110 -344
rect -52 -366 -12 -344
rect 46 -366 86 -344
rect 144 -366 184 -344
rect 242 -366 282 -344
rect 340 -366 380 -344
rect 438 -366 478 -344
rect 536 -366 576 -344
rect 634 -366 674 -344
rect 732 -366 772 -344
rect 830 -366 870 -344
rect 928 -366 968 -344
rect 1026 -366 1066 -344
rect 1124 -366 1164 -344
rect 1222 -366 1262 -344
rect -1130 -788 -1090 -766
rect -1032 -788 -992 -766
rect -934 -788 -894 -766
rect -836 -788 -796 -766
rect -738 -788 -698 -766
rect -640 -788 -600 -766
rect -542 -788 -502 -766
rect -444 -788 -404 -766
rect -346 -788 -306 -766
rect -248 -788 -208 -766
rect -150 -788 -110 -766
rect -52 -788 -12 -766
rect 46 -788 86 -766
rect 144 -788 184 -766
rect 242 -788 282 -766
rect 340 -788 380 -766
rect 438 -788 478 -766
rect 536 -788 576 -766
rect 634 -788 674 -766
rect 732 -788 772 -766
rect 830 -788 870 -766
rect 928 -788 968 -766
rect 1026 -788 1066 -766
rect 1124 -788 1164 -766
rect 1222 -788 1262 -766
rect -1144 -804 1274 -788
rect -1144 -838 -1128 -804
rect -1094 -838 -1029 -804
rect -995 -838 -932 -804
rect -898 -838 -833 -804
rect -799 -838 -736 -804
rect -702 -838 -637 -804
rect -603 -838 -540 -804
rect -506 -838 -441 -804
rect -407 -838 -344 -804
rect -310 -838 -245 -804
rect -211 -838 -148 -804
rect -114 -838 -49 -804
rect -15 -838 48 -804
rect 82 -838 147 -804
rect 181 -838 244 -804
rect 278 -838 343 -804
rect 377 -838 440 -804
rect 474 -838 539 -804
rect 573 -838 636 -804
rect 670 -838 735 -804
rect 769 -838 832 -804
rect 866 -838 931 -804
rect 965 -838 1028 -804
rect 1062 -838 1127 -804
rect 1161 -838 1224 -804
rect 1258 -838 1274 -804
rect -1144 -854 1274 -838
rect -1143 -912 1275 -896
rect -1143 -946 -1127 -912
rect -1093 -946 -1029 -912
rect -995 -946 -931 -912
rect -897 -946 -833 -912
rect -799 -946 -735 -912
rect -701 -946 -637 -912
rect -603 -946 -539 -912
rect -505 -946 -441 -912
rect -407 -946 -343 -912
rect -309 -946 -245 -912
rect -211 -946 -147 -912
rect -113 -946 -49 -912
rect -15 -946 49 -912
rect 83 -946 147 -912
rect 181 -946 245 -912
rect 279 -946 343 -912
rect 377 -946 441 -912
rect 475 -946 539 -912
rect 573 -946 637 -912
rect 671 -946 735 -912
rect 769 -946 833 -912
rect 867 -946 931 -912
rect 965 -946 1029 -912
rect 1063 -946 1127 -912
rect 1161 -946 1225 -912
rect 1259 -946 1275 -912
rect -1143 -962 1275 -946
rect -1130 -984 -1090 -962
rect -1032 -984 -992 -962
rect -934 -984 -894 -962
rect -836 -984 -796 -962
rect -738 -984 -698 -962
rect -640 -984 -600 -962
rect -542 -984 -502 -962
rect -444 -984 -404 -962
rect -346 -984 -306 -962
rect -248 -984 -208 -962
rect -150 -984 -110 -962
rect -52 -984 -12 -962
rect 46 -984 86 -962
rect 144 -984 184 -962
rect 242 -984 282 -962
rect 340 -984 380 -962
rect 438 -984 478 -962
rect 536 -984 576 -962
rect 634 -984 674 -962
rect 732 -984 772 -962
rect 830 -984 870 -962
rect 928 -984 968 -962
rect 1026 -984 1066 -962
rect 1124 -984 1164 -962
rect 1222 -984 1262 -962
rect -1130 -1406 -1090 -1384
rect -1032 -1406 -992 -1384
rect -934 -1406 -894 -1384
rect -836 -1406 -796 -1384
rect -738 -1406 -698 -1384
rect -640 -1406 -600 -1384
rect -542 -1406 -502 -1384
rect -444 -1406 -404 -1384
rect -346 -1406 -306 -1384
rect -248 -1406 -208 -1384
rect -150 -1406 -110 -1384
rect -52 -1406 -12 -1384
rect 46 -1406 86 -1384
rect 144 -1406 184 -1384
rect 242 -1406 282 -1384
rect 340 -1406 380 -1384
rect 438 -1406 478 -1384
rect 536 -1406 576 -1384
rect 634 -1406 674 -1384
rect 732 -1406 772 -1384
rect 830 -1406 870 -1384
rect 928 -1406 968 -1384
rect 1026 -1406 1066 -1384
rect 1124 -1406 1164 -1384
rect 1222 -1406 1262 -1384
rect -1143 -1422 1275 -1406
rect -1143 -1456 -1127 -1422
rect -1093 -1456 -1029 -1422
rect -995 -1456 -931 -1422
rect -897 -1456 -833 -1422
rect -799 -1456 -735 -1422
rect -701 -1456 -637 -1422
rect -603 -1456 -539 -1422
rect -505 -1456 -441 -1422
rect -407 -1456 -343 -1422
rect -309 -1456 -245 -1422
rect -211 -1456 -147 -1422
rect -113 -1456 -49 -1422
rect -15 -1456 49 -1422
rect 83 -1456 147 -1422
rect 181 -1456 245 -1422
rect 279 -1456 343 -1422
rect 377 -1456 441 -1422
rect 475 -1456 539 -1422
rect 573 -1456 637 -1422
rect 671 -1456 735 -1422
rect 769 -1456 833 -1422
rect 867 -1456 931 -1422
rect 965 -1456 1029 -1422
rect 1063 -1456 1127 -1422
rect 1161 -1456 1225 -1422
rect 1259 -1456 1275 -1422
rect -1143 -1472 1275 -1456
rect 2517 830 3955 846
rect 2517 796 2533 830
rect 2567 796 2631 830
rect 2665 796 2729 830
rect 2763 796 2827 830
rect 2861 796 2925 830
rect 2959 796 3023 830
rect 3057 796 3121 830
rect 3155 796 3219 830
rect 3253 796 3317 830
rect 3351 796 3415 830
rect 3449 796 3513 830
rect 3547 796 3611 830
rect 3645 796 3709 830
rect 3743 796 3807 830
rect 3841 796 3905 830
rect 3939 796 3955 830
rect 2517 780 3955 796
rect 2530 758 2570 780
rect 2628 758 2668 780
rect 2726 758 2766 780
rect 2824 758 2864 780
rect 2922 758 2962 780
rect 3020 758 3060 780
rect 3118 758 3158 780
rect 3216 758 3256 780
rect 3314 758 3354 780
rect 3412 758 3452 780
rect 3510 758 3550 780
rect 3608 758 3648 780
rect 3706 758 3746 780
rect 3804 758 3844 780
rect 3902 758 3942 780
rect 2530 336 2570 358
rect 2628 336 2668 358
rect 2726 336 2766 358
rect 2824 336 2864 358
rect 2922 336 2962 358
rect 3020 336 3060 358
rect 3118 336 3158 358
rect 3216 336 3256 358
rect 3314 336 3354 358
rect 3412 336 3452 358
rect 3510 336 3550 358
rect 3608 336 3648 358
rect 3706 336 3746 358
rect 3804 336 3844 358
rect 3902 336 3942 358
rect 2517 320 3955 336
rect 2517 286 2533 320
rect 2567 286 2631 320
rect 2665 286 2729 320
rect 2763 286 2827 320
rect 2861 286 2925 320
rect 2959 286 3023 320
rect 3057 286 3121 320
rect 3155 286 3219 320
rect 3253 286 3317 320
rect 3351 286 3415 320
rect 3449 286 3513 320
rect 3547 286 3611 320
rect 3645 286 3709 320
rect 3743 286 3807 320
rect 3841 286 3905 320
rect 3939 286 3955 320
rect 2517 270 3955 286
rect 2517 212 3955 228
rect 2517 178 2533 212
rect 2567 178 2631 212
rect 2665 178 2729 212
rect 2763 178 2827 212
rect 2861 178 2925 212
rect 2959 178 3023 212
rect 3057 178 3121 212
rect 3155 178 3219 212
rect 3253 178 3317 212
rect 3351 178 3415 212
rect 3449 178 3513 212
rect 3547 178 3611 212
rect 3645 178 3709 212
rect 3743 178 3807 212
rect 3841 178 3905 212
rect 3939 178 3955 212
rect 2517 162 3955 178
rect 2530 140 2570 162
rect 2628 140 2668 162
rect 2726 140 2766 162
rect 2824 140 2864 162
rect 2922 140 2962 162
rect 3020 140 3060 162
rect 3118 140 3158 162
rect 3216 140 3256 162
rect 3314 140 3354 162
rect 3412 140 3452 162
rect 3510 140 3550 162
rect 3608 140 3648 162
rect 3706 140 3746 162
rect 3804 140 3844 162
rect 3902 140 3942 162
rect 2530 -282 2570 -260
rect 2628 -282 2668 -260
rect 2726 -282 2766 -260
rect 2824 -282 2864 -260
rect 2922 -282 2962 -260
rect 3020 -282 3060 -260
rect 3118 -282 3158 -260
rect 3216 -282 3256 -260
rect 3314 -282 3354 -260
rect 3412 -282 3452 -260
rect 3510 -282 3550 -260
rect 3608 -282 3648 -260
rect 3706 -282 3746 -260
rect 3804 -282 3844 -260
rect 3902 -282 3942 -260
rect 2517 -298 3955 -282
rect 2517 -332 2533 -298
rect 2567 -332 2631 -298
rect 2665 -332 2729 -298
rect 2763 -332 2827 -298
rect 2861 -332 2925 -298
rect 2959 -332 3023 -298
rect 3057 -332 3121 -298
rect 3155 -332 3219 -298
rect 3253 -332 3317 -298
rect 3351 -332 3415 -298
rect 3449 -332 3513 -298
rect 3547 -332 3611 -298
rect 3645 -332 3709 -298
rect 3743 -332 3807 -298
rect 3841 -332 3905 -298
rect 3939 -332 3955 -298
rect 2517 -348 3955 -332
rect 1646 -948 2768 -932
rect 1646 -982 1662 -948
rect 1696 -982 1758 -948
rect 1792 -982 1854 -948
rect 1888 -982 1950 -948
rect 1984 -982 2046 -948
rect 2080 -982 2142 -948
rect 2176 -982 2238 -948
rect 2272 -982 2334 -948
rect 2368 -982 2430 -948
rect 2464 -982 2526 -948
rect 2560 -982 2622 -948
rect 2656 -982 2718 -948
rect 2752 -982 2768 -948
rect 1646 -998 2768 -982
rect 1664 -1020 1694 -998
rect 1760 -1020 1790 -998
rect 1856 -1020 1886 -998
rect 1952 -1020 1982 -998
rect 2048 -1020 2078 -998
rect 2144 -1020 2174 -998
rect 2240 -1020 2270 -998
rect 2336 -1020 2366 -998
rect 2432 -1020 2462 -998
rect 2528 -1020 2558 -998
rect 2624 -1020 2654 -998
rect 2720 -1020 2750 -998
rect 1664 -1442 1694 -1420
rect 1760 -1442 1790 -1420
rect 1856 -1442 1886 -1420
rect 1952 -1442 1982 -1420
rect 2048 -1442 2078 -1420
rect 2144 -1442 2174 -1420
rect 2240 -1442 2270 -1420
rect 2336 -1442 2366 -1420
rect 2432 -1442 2462 -1420
rect 2528 -1442 2558 -1420
rect 2624 -1442 2654 -1420
rect 2720 -1442 2750 -1420
rect 1646 -1458 2768 -1442
rect 1646 -1492 1662 -1458
rect 1696 -1492 1758 -1458
rect 1792 -1492 1854 -1458
rect 1888 -1492 1950 -1458
rect 1984 -1492 2046 -1458
rect 2080 -1492 2142 -1458
rect 2176 -1492 2238 -1458
rect 2272 -1492 2334 -1458
rect 2368 -1492 2430 -1458
rect 2464 -1492 2526 -1458
rect 2560 -1492 2622 -1458
rect 2656 -1492 2718 -1458
rect 2752 -1492 2768 -1458
rect 1646 -1508 2768 -1492
rect -1164 -1714 -1098 -1698
rect -1164 -1748 -1148 -1714
rect -1114 -1748 -1098 -1714
rect -1164 -1764 -1098 -1748
rect -972 -1714 -906 -1698
rect -972 -1748 -956 -1714
rect -922 -1748 -906 -1714
rect -1146 -1786 -1116 -1764
rect -1050 -1786 -1020 -1760
rect -972 -1764 -906 -1748
rect -780 -1714 -714 -1698
rect -780 -1748 -764 -1714
rect -730 -1748 -714 -1714
rect -954 -1786 -924 -1764
rect -858 -1786 -828 -1760
rect -780 -1764 -714 -1748
rect -588 -1714 -522 -1698
rect -588 -1748 -572 -1714
rect -538 -1748 -522 -1714
rect -762 -1786 -732 -1764
rect -666 -1786 -636 -1760
rect -588 -1764 -522 -1748
rect -396 -1714 -330 -1698
rect -396 -1748 -380 -1714
rect -346 -1748 -330 -1714
rect -570 -1786 -540 -1764
rect -474 -1786 -444 -1760
rect -396 -1764 -330 -1748
rect -204 -1714 -138 -1698
rect -204 -1748 -188 -1714
rect -154 -1748 -138 -1714
rect -378 -1786 -348 -1764
rect -282 -1786 -252 -1760
rect -204 -1764 -138 -1748
rect -12 -1714 54 -1698
rect -12 -1748 4 -1714
rect 38 -1748 54 -1714
rect -186 -1786 -156 -1764
rect -90 -1786 -60 -1760
rect -12 -1764 54 -1748
rect 180 -1714 246 -1698
rect 180 -1748 196 -1714
rect 230 -1748 246 -1714
rect 6 -1786 36 -1764
rect 102 -1786 132 -1760
rect 180 -1764 246 -1748
rect 372 -1714 438 -1698
rect 372 -1748 388 -1714
rect 422 -1748 438 -1714
rect 198 -1786 228 -1764
rect 294 -1786 324 -1760
rect 372 -1764 438 -1748
rect 564 -1714 630 -1698
rect 564 -1748 580 -1714
rect 614 -1748 630 -1714
rect 390 -1786 420 -1764
rect 486 -1786 516 -1760
rect 564 -1764 630 -1748
rect 756 -1714 822 -1698
rect 756 -1748 772 -1714
rect 806 -1748 822 -1714
rect 582 -1786 612 -1764
rect 678 -1786 708 -1760
rect 756 -1764 822 -1748
rect 948 -1714 1014 -1698
rect 948 -1748 964 -1714
rect 998 -1748 1014 -1714
rect 774 -1786 804 -1764
rect 870 -1786 900 -1760
rect 948 -1764 1014 -1748
rect 1140 -1714 1206 -1698
rect 1140 -1748 1156 -1714
rect 1190 -1748 1206 -1714
rect 966 -1786 996 -1764
rect 1062 -1786 1092 -1760
rect 1140 -1764 1206 -1748
rect 1158 -1786 1188 -1764
rect -1146 -2212 -1116 -2186
rect -1050 -2208 -1020 -2186
rect -1068 -2224 -1002 -2208
rect -954 -2212 -924 -2186
rect -858 -2208 -828 -2186
rect -1068 -2258 -1052 -2224
rect -1018 -2258 -1002 -2224
rect -1068 -2274 -1002 -2258
rect -876 -2224 -810 -2208
rect -762 -2212 -732 -2186
rect -666 -2208 -636 -2186
rect -876 -2258 -860 -2224
rect -826 -2258 -810 -2224
rect -876 -2274 -810 -2258
rect -684 -2224 -618 -2208
rect -570 -2212 -540 -2186
rect -474 -2208 -444 -2186
rect -684 -2258 -668 -2224
rect -634 -2258 -618 -2224
rect -684 -2274 -618 -2258
rect -492 -2224 -426 -2208
rect -378 -2212 -348 -2186
rect -282 -2208 -252 -2186
rect -492 -2258 -476 -2224
rect -442 -2258 -426 -2224
rect -492 -2274 -426 -2258
rect -300 -2224 -234 -2208
rect -186 -2212 -156 -2186
rect -90 -2208 -60 -2186
rect -300 -2258 -284 -2224
rect -250 -2258 -234 -2224
rect -300 -2274 -234 -2258
rect -108 -2224 -42 -2208
rect 6 -2212 36 -2186
rect 102 -2208 132 -2186
rect -108 -2258 -92 -2224
rect -58 -2258 -42 -2224
rect -108 -2274 -42 -2258
rect 84 -2224 150 -2208
rect 198 -2212 228 -2186
rect 294 -2208 324 -2186
rect 84 -2258 100 -2224
rect 134 -2258 150 -2224
rect 84 -2274 150 -2258
rect 276 -2224 342 -2208
rect 390 -2212 420 -2186
rect 486 -2208 516 -2186
rect 276 -2258 292 -2224
rect 326 -2258 342 -2224
rect 276 -2274 342 -2258
rect 468 -2224 534 -2208
rect 582 -2212 612 -2186
rect 678 -2208 708 -2186
rect 468 -2258 484 -2224
rect 518 -2258 534 -2224
rect 468 -2274 534 -2258
rect 660 -2224 726 -2208
rect 774 -2212 804 -2186
rect 870 -2208 900 -2186
rect 660 -2258 676 -2224
rect 710 -2258 726 -2224
rect 660 -2274 726 -2258
rect 852 -2224 918 -2208
rect 966 -2212 996 -2186
rect 1062 -2208 1092 -2186
rect 852 -2258 868 -2224
rect 902 -2258 918 -2224
rect 852 -2274 918 -2258
rect 1044 -2224 1110 -2208
rect 1158 -2212 1188 -2186
rect 1044 -2258 1060 -2224
rect 1094 -2258 1110 -2224
rect 1044 -2274 1110 -2258
rect -1068 -2332 -1002 -2316
rect -1068 -2366 -1052 -2332
rect -1018 -2366 -1002 -2332
rect -1146 -2404 -1116 -2378
rect -1068 -2382 -1002 -2366
rect -876 -2332 -810 -2316
rect -876 -2366 -860 -2332
rect -826 -2366 -810 -2332
rect -1050 -2404 -1020 -2382
rect -954 -2404 -924 -2378
rect -876 -2382 -810 -2366
rect -684 -2332 -618 -2316
rect -684 -2366 -668 -2332
rect -634 -2366 -618 -2332
rect -858 -2404 -828 -2382
rect -762 -2404 -732 -2378
rect -684 -2382 -618 -2366
rect -492 -2332 -426 -2316
rect -492 -2366 -476 -2332
rect -442 -2366 -426 -2332
rect -666 -2404 -636 -2382
rect -570 -2404 -540 -2378
rect -492 -2382 -426 -2366
rect -300 -2332 -234 -2316
rect -300 -2366 -284 -2332
rect -250 -2366 -234 -2332
rect -474 -2404 -444 -2382
rect -378 -2404 -348 -2378
rect -300 -2382 -234 -2366
rect -108 -2332 -42 -2316
rect -108 -2366 -92 -2332
rect -58 -2366 -42 -2332
rect -282 -2404 -252 -2382
rect -186 -2404 -156 -2378
rect -108 -2382 -42 -2366
rect 84 -2332 150 -2316
rect 84 -2366 100 -2332
rect 134 -2366 150 -2332
rect -90 -2404 -60 -2382
rect 6 -2404 36 -2378
rect 84 -2382 150 -2366
rect 276 -2332 342 -2316
rect 276 -2366 292 -2332
rect 326 -2366 342 -2332
rect 102 -2404 132 -2382
rect 198 -2404 228 -2378
rect 276 -2382 342 -2366
rect 468 -2332 534 -2316
rect 468 -2366 484 -2332
rect 518 -2366 534 -2332
rect 294 -2404 324 -2382
rect 390 -2404 420 -2378
rect 468 -2382 534 -2366
rect 660 -2332 726 -2316
rect 660 -2366 676 -2332
rect 710 -2366 726 -2332
rect 486 -2404 516 -2382
rect 582 -2404 612 -2378
rect 660 -2382 726 -2366
rect 852 -2332 918 -2316
rect 852 -2366 868 -2332
rect 902 -2366 918 -2332
rect 678 -2404 708 -2382
rect 774 -2404 804 -2378
rect 852 -2382 918 -2366
rect 1044 -2332 1110 -2316
rect 1044 -2366 1060 -2332
rect 1094 -2366 1110 -2332
rect 870 -2404 900 -2382
rect 966 -2404 996 -2378
rect 1044 -2382 1110 -2366
rect 1062 -2404 1092 -2382
rect 1158 -2404 1188 -2378
rect -1146 -2826 -1116 -2804
rect -1164 -2842 -1098 -2826
rect -1050 -2830 -1020 -2804
rect -954 -2826 -924 -2804
rect -1164 -2876 -1148 -2842
rect -1114 -2876 -1098 -2842
rect -1164 -2892 -1098 -2876
rect -972 -2842 -906 -2826
rect -858 -2830 -828 -2804
rect -762 -2826 -732 -2804
rect -972 -2876 -956 -2842
rect -922 -2876 -906 -2842
rect -972 -2892 -906 -2876
rect -780 -2842 -714 -2826
rect -666 -2830 -636 -2804
rect -570 -2826 -540 -2804
rect -780 -2876 -764 -2842
rect -730 -2876 -714 -2842
rect -780 -2892 -714 -2876
rect -588 -2842 -522 -2826
rect -474 -2830 -444 -2804
rect -378 -2826 -348 -2804
rect -588 -2876 -572 -2842
rect -538 -2876 -522 -2842
rect -588 -2892 -522 -2876
rect -396 -2842 -330 -2826
rect -282 -2830 -252 -2804
rect -186 -2826 -156 -2804
rect -396 -2876 -380 -2842
rect -346 -2876 -330 -2842
rect -396 -2892 -330 -2876
rect -204 -2842 -138 -2826
rect -90 -2830 -60 -2804
rect 6 -2826 36 -2804
rect -204 -2876 -188 -2842
rect -154 -2876 -138 -2842
rect -204 -2892 -138 -2876
rect -12 -2842 54 -2826
rect 102 -2830 132 -2804
rect 198 -2826 228 -2804
rect -12 -2876 4 -2842
rect 38 -2876 54 -2842
rect -12 -2892 54 -2876
rect 180 -2842 246 -2826
rect 294 -2830 324 -2804
rect 390 -2826 420 -2804
rect 180 -2876 196 -2842
rect 230 -2876 246 -2842
rect 180 -2892 246 -2876
rect 372 -2842 438 -2826
rect 486 -2830 516 -2804
rect 582 -2826 612 -2804
rect 372 -2876 388 -2842
rect 422 -2876 438 -2842
rect 372 -2892 438 -2876
rect 564 -2842 630 -2826
rect 678 -2830 708 -2804
rect 774 -2826 804 -2804
rect 564 -2876 580 -2842
rect 614 -2876 630 -2842
rect 564 -2892 630 -2876
rect 756 -2842 822 -2826
rect 870 -2830 900 -2804
rect 966 -2826 996 -2804
rect 756 -2876 772 -2842
rect 806 -2876 822 -2842
rect 756 -2892 822 -2876
rect 948 -2842 1014 -2826
rect 1062 -2830 1092 -2804
rect 1158 -2826 1188 -2804
rect 948 -2876 964 -2842
rect 998 -2876 1014 -2842
rect 948 -2892 1014 -2876
rect 1140 -2842 1206 -2826
rect 1140 -2876 1156 -2842
rect 1190 -2876 1206 -2842
rect 1140 -2892 1206 -2876
rect -1164 -2950 -1098 -2934
rect -1164 -2984 -1148 -2950
rect -1114 -2984 -1098 -2950
rect -1164 -3000 -1098 -2984
rect -972 -2950 -906 -2934
rect -972 -2984 -956 -2950
rect -922 -2984 -906 -2950
rect -1146 -3022 -1116 -3000
rect -1050 -3022 -1020 -2996
rect -972 -3000 -906 -2984
rect -780 -2950 -714 -2934
rect -780 -2984 -764 -2950
rect -730 -2984 -714 -2950
rect -954 -3022 -924 -3000
rect -858 -3022 -828 -2996
rect -780 -3000 -714 -2984
rect -588 -2950 -522 -2934
rect -588 -2984 -572 -2950
rect -538 -2984 -522 -2950
rect -762 -3022 -732 -3000
rect -666 -3022 -636 -2996
rect -588 -3000 -522 -2984
rect -396 -2950 -330 -2934
rect -396 -2984 -380 -2950
rect -346 -2984 -330 -2950
rect -570 -3022 -540 -3000
rect -474 -3022 -444 -2996
rect -396 -3000 -330 -2984
rect -204 -2950 -138 -2934
rect -204 -2984 -188 -2950
rect -154 -2984 -138 -2950
rect -378 -3022 -348 -3000
rect -282 -3022 -252 -2996
rect -204 -3000 -138 -2984
rect -12 -2950 54 -2934
rect -12 -2984 4 -2950
rect 38 -2984 54 -2950
rect -186 -3022 -156 -3000
rect -90 -3022 -60 -2996
rect -12 -3000 54 -2984
rect 180 -2950 246 -2934
rect 180 -2984 196 -2950
rect 230 -2984 246 -2950
rect 6 -3022 36 -3000
rect 102 -3022 132 -2996
rect 180 -3000 246 -2984
rect 372 -2950 438 -2934
rect 372 -2984 388 -2950
rect 422 -2984 438 -2950
rect 198 -3022 228 -3000
rect 294 -3022 324 -2996
rect 372 -3000 438 -2984
rect 564 -2950 630 -2934
rect 564 -2984 580 -2950
rect 614 -2984 630 -2950
rect 390 -3022 420 -3000
rect 486 -3022 516 -2996
rect 564 -3000 630 -2984
rect 756 -2950 822 -2934
rect 756 -2984 772 -2950
rect 806 -2984 822 -2950
rect 582 -3022 612 -3000
rect 678 -3022 708 -2996
rect 756 -3000 822 -2984
rect 948 -2950 1014 -2934
rect 948 -2984 964 -2950
rect 998 -2984 1014 -2950
rect 774 -3022 804 -3000
rect 870 -3022 900 -2996
rect 948 -3000 1014 -2984
rect 1140 -2950 1206 -2934
rect 1140 -2984 1156 -2950
rect 1190 -2984 1206 -2950
rect 966 -3022 996 -3000
rect 1062 -3022 1092 -2996
rect 1140 -3000 1206 -2984
rect 1158 -3022 1188 -3000
rect -1146 -3448 -1116 -3422
rect -1050 -3444 -1020 -3422
rect -1068 -3460 -1002 -3444
rect -954 -3448 -924 -3422
rect -858 -3444 -828 -3422
rect -1068 -3494 -1052 -3460
rect -1018 -3494 -1002 -3460
rect -1068 -3510 -1002 -3494
rect -876 -3460 -810 -3444
rect -762 -3448 -732 -3422
rect -666 -3444 -636 -3422
rect -876 -3494 -860 -3460
rect -826 -3494 -810 -3460
rect -876 -3510 -810 -3494
rect -684 -3460 -618 -3444
rect -570 -3448 -540 -3422
rect -474 -3444 -444 -3422
rect -684 -3494 -668 -3460
rect -634 -3494 -618 -3460
rect -684 -3510 -618 -3494
rect -492 -3460 -426 -3444
rect -378 -3448 -348 -3422
rect -282 -3444 -252 -3422
rect -492 -3494 -476 -3460
rect -442 -3494 -426 -3460
rect -492 -3510 -426 -3494
rect -300 -3460 -234 -3444
rect -186 -3448 -156 -3422
rect -90 -3444 -60 -3422
rect -300 -3494 -284 -3460
rect -250 -3494 -234 -3460
rect -300 -3510 -234 -3494
rect -108 -3460 -42 -3444
rect 6 -3448 36 -3422
rect 102 -3444 132 -3422
rect -108 -3494 -92 -3460
rect -58 -3494 -42 -3460
rect -108 -3510 -42 -3494
rect 84 -3460 150 -3444
rect 198 -3448 228 -3422
rect 294 -3444 324 -3422
rect 84 -3494 100 -3460
rect 134 -3494 150 -3460
rect 84 -3510 150 -3494
rect 276 -3460 342 -3444
rect 390 -3448 420 -3422
rect 486 -3444 516 -3422
rect 276 -3494 292 -3460
rect 326 -3494 342 -3460
rect 276 -3510 342 -3494
rect 468 -3460 534 -3444
rect 582 -3448 612 -3422
rect 678 -3444 708 -3422
rect 468 -3494 484 -3460
rect 518 -3494 534 -3460
rect 468 -3510 534 -3494
rect 660 -3460 726 -3444
rect 774 -3448 804 -3422
rect 870 -3444 900 -3422
rect 660 -3494 676 -3460
rect 710 -3494 726 -3460
rect 660 -3510 726 -3494
rect 852 -3460 918 -3444
rect 966 -3448 996 -3422
rect 1062 -3444 1092 -3422
rect 852 -3494 868 -3460
rect 902 -3494 918 -3460
rect 852 -3510 918 -3494
rect 1044 -3460 1110 -3444
rect 1158 -3448 1188 -3422
rect 1044 -3494 1060 -3460
rect 1094 -3494 1110 -3460
rect 1044 -3510 1110 -3494
rect -1068 -3568 -1002 -3552
rect -1068 -3602 -1052 -3568
rect -1018 -3602 -1002 -3568
rect -1146 -3640 -1116 -3614
rect -1068 -3618 -1002 -3602
rect -876 -3568 -810 -3552
rect -876 -3602 -860 -3568
rect -826 -3602 -810 -3568
rect -1050 -3640 -1020 -3618
rect -954 -3640 -924 -3614
rect -876 -3618 -810 -3602
rect -684 -3568 -618 -3552
rect -684 -3602 -668 -3568
rect -634 -3602 -618 -3568
rect -858 -3640 -828 -3618
rect -762 -3640 -732 -3614
rect -684 -3618 -618 -3602
rect -492 -3568 -426 -3552
rect -492 -3602 -476 -3568
rect -442 -3602 -426 -3568
rect -666 -3640 -636 -3618
rect -570 -3640 -540 -3614
rect -492 -3618 -426 -3602
rect -300 -3568 -234 -3552
rect -300 -3602 -284 -3568
rect -250 -3602 -234 -3568
rect -474 -3640 -444 -3618
rect -378 -3640 -348 -3614
rect -300 -3618 -234 -3602
rect -108 -3568 -42 -3552
rect -108 -3602 -92 -3568
rect -58 -3602 -42 -3568
rect -282 -3640 -252 -3618
rect -186 -3640 -156 -3614
rect -108 -3618 -42 -3602
rect 84 -3568 150 -3552
rect 84 -3602 100 -3568
rect 134 -3602 150 -3568
rect -90 -3640 -60 -3618
rect 6 -3640 36 -3614
rect 84 -3618 150 -3602
rect 276 -3568 342 -3552
rect 276 -3602 292 -3568
rect 326 -3602 342 -3568
rect 102 -3640 132 -3618
rect 198 -3640 228 -3614
rect 276 -3618 342 -3602
rect 468 -3568 534 -3552
rect 468 -3602 484 -3568
rect 518 -3602 534 -3568
rect 294 -3640 324 -3618
rect 390 -3640 420 -3614
rect 468 -3618 534 -3602
rect 660 -3568 726 -3552
rect 660 -3602 676 -3568
rect 710 -3602 726 -3568
rect 486 -3640 516 -3618
rect 582 -3640 612 -3614
rect 660 -3618 726 -3602
rect 852 -3568 918 -3552
rect 852 -3602 868 -3568
rect 902 -3602 918 -3568
rect 678 -3640 708 -3618
rect 774 -3640 804 -3614
rect 852 -3618 918 -3602
rect 1044 -3568 1110 -3552
rect 1044 -3602 1060 -3568
rect 1094 -3602 1110 -3568
rect 870 -3640 900 -3618
rect 966 -3640 996 -3614
rect 1044 -3618 1110 -3602
rect 1062 -3640 1092 -3618
rect 1158 -3640 1188 -3614
rect -1146 -4062 -1116 -4040
rect -1164 -4078 -1098 -4062
rect -1050 -4066 -1020 -4040
rect -954 -4062 -924 -4040
rect -1164 -4112 -1148 -4078
rect -1114 -4112 -1098 -4078
rect -1164 -4128 -1098 -4112
rect -972 -4078 -906 -4062
rect -858 -4066 -828 -4040
rect -762 -4062 -732 -4040
rect -972 -4112 -956 -4078
rect -922 -4112 -906 -4078
rect -972 -4128 -906 -4112
rect -780 -4078 -714 -4062
rect -666 -4066 -636 -4040
rect -570 -4062 -540 -4040
rect -780 -4112 -764 -4078
rect -730 -4112 -714 -4078
rect -780 -4128 -714 -4112
rect -588 -4078 -522 -4062
rect -474 -4066 -444 -4040
rect -378 -4062 -348 -4040
rect -588 -4112 -572 -4078
rect -538 -4112 -522 -4078
rect -588 -4128 -522 -4112
rect -396 -4078 -330 -4062
rect -282 -4066 -252 -4040
rect -186 -4062 -156 -4040
rect -396 -4112 -380 -4078
rect -346 -4112 -330 -4078
rect -396 -4128 -330 -4112
rect -204 -4078 -138 -4062
rect -90 -4066 -60 -4040
rect 6 -4062 36 -4040
rect -204 -4112 -188 -4078
rect -154 -4112 -138 -4078
rect -204 -4128 -138 -4112
rect -12 -4078 54 -4062
rect 102 -4066 132 -4040
rect 198 -4062 228 -4040
rect -12 -4112 4 -4078
rect 38 -4112 54 -4078
rect -12 -4128 54 -4112
rect 180 -4078 246 -4062
rect 294 -4066 324 -4040
rect 390 -4062 420 -4040
rect 180 -4112 196 -4078
rect 230 -4112 246 -4078
rect 180 -4128 246 -4112
rect 372 -4078 438 -4062
rect 486 -4066 516 -4040
rect 582 -4062 612 -4040
rect 372 -4112 388 -4078
rect 422 -4112 438 -4078
rect 372 -4128 438 -4112
rect 564 -4078 630 -4062
rect 678 -4066 708 -4040
rect 774 -4062 804 -4040
rect 564 -4112 580 -4078
rect 614 -4112 630 -4078
rect 564 -4128 630 -4112
rect 756 -4078 822 -4062
rect 870 -4066 900 -4040
rect 966 -4062 996 -4040
rect 756 -4112 772 -4078
rect 806 -4112 822 -4078
rect 756 -4128 822 -4112
rect 948 -4078 1014 -4062
rect 1062 -4066 1092 -4040
rect 1158 -4062 1188 -4040
rect 948 -4112 964 -4078
rect 998 -4112 1014 -4078
rect 948 -4128 1014 -4112
rect 1140 -4078 1206 -4062
rect 1140 -4112 1156 -4078
rect 1190 -4112 1206 -4078
rect 1140 -4128 1206 -4112
rect 1660 -1768 1860 -1752
rect 1660 -1802 1676 -1768
rect 1844 -1802 1860 -1768
rect 1660 -1840 1860 -1802
rect 1918 -1768 2118 -1752
rect 1918 -1802 1934 -1768
rect 2102 -1802 2118 -1768
rect 1918 -1840 2118 -1802
rect 2176 -1768 2376 -1752
rect 2176 -1802 2192 -1768
rect 2360 -1802 2376 -1768
rect 2176 -1840 2376 -1802
rect 2434 -1768 2634 -1752
rect 2434 -1802 2450 -1768
rect 2618 -1802 2634 -1768
rect 2434 -1840 2634 -1802
rect 2692 -1768 2892 -1752
rect 2692 -1802 2708 -1768
rect 2876 -1802 2892 -1768
rect 2692 -1840 2892 -1802
rect 2950 -1768 3150 -1752
rect 2950 -1802 2966 -1768
rect 3134 -1802 3150 -1768
rect 2950 -1840 3150 -1802
rect 1660 -2278 1860 -2240
rect 1660 -2312 1676 -2278
rect 1844 -2312 1860 -2278
rect 1660 -2328 1860 -2312
rect 1918 -2278 2118 -2240
rect 1918 -2312 1934 -2278
rect 2102 -2312 2118 -2278
rect 1918 -2328 2118 -2312
rect 2176 -2278 2376 -2240
rect 2176 -2312 2192 -2278
rect 2360 -2312 2376 -2278
rect 2176 -2328 2376 -2312
rect 2434 -2278 2634 -2240
rect 2434 -2312 2450 -2278
rect 2618 -2312 2634 -2278
rect 2434 -2328 2634 -2312
rect 2692 -2278 2892 -2240
rect 2692 -2312 2708 -2278
rect 2876 -2312 2892 -2278
rect 2692 -2328 2892 -2312
rect 2950 -2278 3150 -2240
rect 2950 -2312 2966 -2278
rect 3134 -2312 3150 -2278
rect 2950 -2328 3150 -2312
rect -1143 -4444 295 -4428
rect -1143 -4478 -1127 -4444
rect -1093 -4478 -1029 -4444
rect -995 -4478 -931 -4444
rect -897 -4478 -833 -4444
rect -799 -4478 -735 -4444
rect -701 -4478 -637 -4444
rect -603 -4478 -539 -4444
rect -505 -4478 -441 -4444
rect -407 -4478 -343 -4444
rect -309 -4478 -245 -4444
rect -211 -4478 -147 -4444
rect -113 -4478 -49 -4444
rect -15 -4478 49 -4444
rect 83 -4478 147 -4444
rect 181 -4478 245 -4444
rect 279 -4478 295 -4444
rect -1143 -4494 295 -4478
rect -1130 -4525 -1090 -4494
rect -1032 -4525 -992 -4494
rect -934 -4525 -894 -4494
rect -836 -4525 -796 -4494
rect -738 -4525 -698 -4494
rect -640 -4525 -600 -4494
rect -542 -4525 -502 -4494
rect -444 -4525 -404 -4494
rect -346 -4525 -306 -4494
rect -248 -4525 -208 -4494
rect -150 -4525 -110 -4494
rect -52 -4525 -12 -4494
rect 46 -4525 86 -4494
rect 144 -4525 184 -4494
rect 242 -4525 282 -4494
rect -1130 -4956 -1090 -4925
rect -1032 -4956 -992 -4925
rect -934 -4956 -894 -4925
rect -836 -4956 -796 -4925
rect -738 -4956 -698 -4925
rect -640 -4956 -600 -4925
rect -542 -4956 -502 -4925
rect -444 -4956 -404 -4925
rect -346 -4956 -306 -4925
rect -248 -4956 -208 -4925
rect -150 -4956 -110 -4925
rect -52 -4956 -12 -4925
rect 46 -4956 86 -4925
rect 144 -4956 184 -4925
rect 242 -4956 282 -4925
rect -1143 -4972 295 -4956
rect -1143 -5006 -1127 -4972
rect -1093 -5006 -1029 -4972
rect -995 -5006 -931 -4972
rect -897 -5006 -833 -4972
rect -799 -5006 -735 -4972
rect -701 -5006 -637 -4972
rect -603 -5006 -539 -4972
rect -505 -5006 -441 -4972
rect -407 -5006 -343 -4972
rect -309 -5006 -245 -4972
rect -211 -5006 -147 -4972
rect -113 -5006 -49 -4972
rect -15 -5006 49 -4972
rect 83 -5006 147 -4972
rect 181 -5006 245 -4972
rect 279 -5006 295 -4972
rect -1143 -5022 295 -5006
rect -1143 -5080 295 -5064
rect -1143 -5114 -1127 -5080
rect -1093 -5114 -1029 -5080
rect -995 -5114 -931 -5080
rect -897 -5114 -833 -5080
rect -799 -5114 -735 -5080
rect -701 -5114 -637 -5080
rect -603 -5114 -539 -5080
rect -505 -5114 -441 -5080
rect -407 -5114 -343 -5080
rect -309 -5114 -245 -5080
rect -211 -5114 -147 -5080
rect -113 -5114 -49 -5080
rect -15 -5114 49 -5080
rect 83 -5114 147 -5080
rect 181 -5114 245 -5080
rect 279 -5114 295 -5080
rect -1143 -5130 295 -5114
rect -1130 -5161 -1090 -5130
rect -1032 -5161 -992 -5130
rect -934 -5161 -894 -5130
rect -836 -5161 -796 -5130
rect -738 -5161 -698 -5130
rect -640 -5161 -600 -5130
rect -542 -5161 -502 -5130
rect -444 -5161 -404 -5130
rect -346 -5161 -306 -5130
rect -248 -5161 -208 -5130
rect -150 -5161 -110 -5130
rect -52 -5161 -12 -5130
rect 46 -5161 86 -5130
rect 144 -5161 184 -5130
rect 242 -5161 282 -5130
rect -1130 -5592 -1090 -5561
rect -1032 -5592 -992 -5561
rect -934 -5592 -894 -5561
rect -836 -5592 -796 -5561
rect -738 -5592 -698 -5561
rect -640 -5592 -600 -5561
rect -542 -5592 -502 -5561
rect -444 -5592 -404 -5561
rect -346 -5592 -306 -5561
rect -248 -5592 -208 -5561
rect -150 -5592 -110 -5561
rect -52 -5592 -12 -5561
rect 46 -5592 86 -5561
rect 144 -5592 184 -5561
rect 242 -5592 282 -5561
rect -1143 -5608 295 -5592
rect -1143 -5642 -1127 -5608
rect -1093 -5642 -1029 -5608
rect -995 -5642 -931 -5608
rect -897 -5642 -833 -5608
rect -799 -5642 -735 -5608
rect -701 -5642 -637 -5608
rect -603 -5642 -539 -5608
rect -505 -5642 -441 -5608
rect -407 -5642 -343 -5608
rect -309 -5642 -245 -5608
rect -211 -5642 -147 -5608
rect -113 -5642 -49 -5608
rect -15 -5642 49 -5608
rect 83 -5642 147 -5608
rect 181 -5642 245 -5608
rect 279 -5642 295 -5608
rect -1143 -5658 295 -5642
rect 655 -4444 2093 -4428
rect 655 -4478 671 -4444
rect 705 -4478 769 -4444
rect 803 -4478 867 -4444
rect 901 -4478 965 -4444
rect 999 -4478 1063 -4444
rect 1097 -4478 1161 -4444
rect 1195 -4478 1259 -4444
rect 1293 -4478 1357 -4444
rect 1391 -4478 1455 -4444
rect 1489 -4478 1553 -4444
rect 1587 -4478 1651 -4444
rect 1685 -4478 1749 -4444
rect 1783 -4478 1847 -4444
rect 1881 -4478 1945 -4444
rect 1979 -4478 2043 -4444
rect 2077 -4478 2093 -4444
rect 655 -4494 2093 -4478
rect 668 -4525 708 -4494
rect 766 -4525 806 -4494
rect 864 -4525 904 -4494
rect 962 -4525 1002 -4494
rect 1060 -4525 1100 -4494
rect 1158 -4525 1198 -4494
rect 1256 -4525 1296 -4494
rect 1354 -4525 1394 -4494
rect 1452 -4525 1492 -4494
rect 1550 -4525 1590 -4494
rect 1648 -4525 1688 -4494
rect 1746 -4525 1786 -4494
rect 1844 -4525 1884 -4494
rect 1942 -4525 1982 -4494
rect 2040 -4525 2080 -4494
rect 668 -4956 708 -4925
rect 766 -4956 806 -4925
rect 864 -4956 904 -4925
rect 962 -4956 1002 -4925
rect 1060 -4956 1100 -4925
rect 1158 -4956 1198 -4925
rect 1256 -4956 1296 -4925
rect 1354 -4956 1394 -4925
rect 1452 -4956 1492 -4925
rect 1550 -4956 1590 -4925
rect 1648 -4956 1688 -4925
rect 1746 -4956 1786 -4925
rect 1844 -4956 1884 -4925
rect 1942 -4956 1982 -4925
rect 2040 -4956 2080 -4925
rect 655 -4972 2093 -4956
rect 655 -5006 671 -4972
rect 705 -5006 769 -4972
rect 803 -5006 867 -4972
rect 901 -5006 965 -4972
rect 999 -5006 1063 -4972
rect 1097 -5006 1161 -4972
rect 1195 -5006 1259 -4972
rect 1293 -5006 1357 -4972
rect 1391 -5006 1455 -4972
rect 1489 -5006 1553 -4972
rect 1587 -5006 1651 -4972
rect 1685 -5006 1749 -4972
rect 1783 -5006 1847 -4972
rect 1881 -5006 1945 -4972
rect 1979 -5006 2043 -4972
rect 2077 -5006 2093 -4972
rect 655 -5022 2093 -5006
rect 655 -5080 2093 -5064
rect 655 -5114 671 -5080
rect 705 -5114 769 -5080
rect 803 -5114 867 -5080
rect 901 -5114 965 -5080
rect 999 -5114 1063 -5080
rect 1097 -5114 1161 -5080
rect 1195 -5114 1259 -5080
rect 1293 -5114 1357 -5080
rect 1391 -5114 1455 -5080
rect 1489 -5114 1553 -5080
rect 1587 -5114 1651 -5080
rect 1685 -5114 1749 -5080
rect 1783 -5114 1847 -5080
rect 1881 -5114 1945 -5080
rect 1979 -5114 2043 -5080
rect 2077 -5114 2093 -5080
rect 655 -5130 2093 -5114
rect 668 -5161 708 -5130
rect 766 -5161 806 -5130
rect 864 -5161 904 -5130
rect 962 -5161 1002 -5130
rect 1060 -5161 1100 -5130
rect 1158 -5161 1198 -5130
rect 1256 -5161 1296 -5130
rect 1354 -5161 1394 -5130
rect 1452 -5161 1492 -5130
rect 1550 -5161 1590 -5130
rect 1648 -5161 1688 -5130
rect 1746 -5161 1786 -5130
rect 1844 -5161 1884 -5130
rect 1942 -5161 1982 -5130
rect 2040 -5161 2080 -5130
rect 668 -5592 708 -5561
rect 766 -5592 806 -5561
rect 864 -5592 904 -5561
rect 962 -5592 1002 -5561
rect 1060 -5592 1100 -5561
rect 1158 -5592 1198 -5561
rect 1256 -5592 1296 -5561
rect 1354 -5592 1394 -5561
rect 1452 -5592 1492 -5561
rect 1550 -5592 1590 -5561
rect 1648 -5592 1688 -5561
rect 1746 -5592 1786 -5561
rect 1844 -5592 1884 -5561
rect 1942 -5592 1982 -5561
rect 2040 -5592 2080 -5561
rect 655 -5608 2093 -5592
rect 655 -5642 671 -5608
rect 705 -5642 769 -5608
rect 803 -5642 867 -5608
rect 901 -5642 965 -5608
rect 999 -5642 1063 -5608
rect 1097 -5642 1161 -5608
rect 1195 -5642 1259 -5608
rect 1293 -5642 1357 -5608
rect 1391 -5642 1455 -5608
rect 1489 -5642 1553 -5608
rect 1587 -5642 1651 -5608
rect 1685 -5642 1749 -5608
rect 1783 -5642 1847 -5608
rect 1881 -5642 1945 -5608
rect 1979 -5642 2043 -5608
rect 2077 -5642 2093 -5608
rect 655 -5658 2093 -5642
rect 2470 -5096 2570 -5080
rect 2470 -5130 2486 -5096
rect 2554 -5130 2570 -5096
rect 2470 -5177 2570 -5130
rect 2628 -5096 2728 -5080
rect 2628 -5130 2644 -5096
rect 2712 -5130 2728 -5096
rect 2628 -5177 2728 -5130
rect 2786 -5096 2886 -5080
rect 2786 -5130 2802 -5096
rect 2870 -5130 2886 -5096
rect 2786 -5177 2886 -5130
rect 2944 -5096 3044 -5080
rect 2944 -5130 2960 -5096
rect 3028 -5130 3044 -5096
rect 2944 -5177 3044 -5130
rect 3102 -5096 3202 -5080
rect 3102 -5130 3118 -5096
rect 3186 -5130 3202 -5096
rect 3102 -5177 3202 -5130
rect 3260 -5096 3360 -5080
rect 3260 -5130 3276 -5096
rect 3344 -5130 3360 -5096
rect 3260 -5177 3360 -5130
rect 3418 -5096 3518 -5080
rect 3418 -5130 3434 -5096
rect 3502 -5130 3518 -5096
rect 3418 -5177 3518 -5130
rect 3576 -5096 3676 -5080
rect 3576 -5130 3592 -5096
rect 3660 -5130 3676 -5096
rect 3576 -5177 3676 -5130
rect 3734 -5096 3834 -5080
rect 3734 -5130 3750 -5096
rect 3818 -5130 3834 -5096
rect 3734 -5177 3834 -5130
rect 3892 -5096 3992 -5080
rect 3892 -5130 3908 -5096
rect 3976 -5130 3992 -5096
rect 3892 -5177 3992 -5130
rect 2470 -5624 2570 -5577
rect 2470 -5658 2486 -5624
rect 2554 -5658 2570 -5624
rect 2470 -5674 2570 -5658
rect 2628 -5624 2728 -5577
rect 2628 -5658 2644 -5624
rect 2712 -5658 2728 -5624
rect 2628 -5674 2728 -5658
rect 2786 -5624 2886 -5577
rect 2786 -5658 2802 -5624
rect 2870 -5658 2886 -5624
rect 2786 -5674 2886 -5658
rect 2944 -5624 3044 -5577
rect 2944 -5658 2960 -5624
rect 3028 -5658 3044 -5624
rect 2944 -5674 3044 -5658
rect 3102 -5624 3202 -5577
rect 3102 -5658 3118 -5624
rect 3186 -5658 3202 -5624
rect 3102 -5674 3202 -5658
rect 3260 -5624 3360 -5577
rect 3260 -5658 3276 -5624
rect 3344 -5658 3360 -5624
rect 3260 -5674 3360 -5658
rect 3418 -5624 3518 -5577
rect 3418 -5658 3434 -5624
rect 3502 -5658 3518 -5624
rect 3418 -5674 3518 -5658
rect 3576 -5624 3676 -5577
rect 3576 -5658 3592 -5624
rect 3660 -5658 3676 -5624
rect 3576 -5674 3676 -5658
rect 3734 -5624 3834 -5577
rect 3734 -5658 3750 -5624
rect 3818 -5658 3834 -5624
rect 3734 -5674 3834 -5658
rect 3892 -5624 3992 -5577
rect 3892 -5658 3908 -5624
rect 3976 -5658 3992 -5624
rect 3892 -5674 3992 -5658
rect -1144 -5920 1275 -5904
rect -1144 -5954 -1127 -5920
rect -1093 -5954 -1030 -5920
rect -996 -5954 -931 -5920
rect -897 -5954 -834 -5920
rect -800 -5954 -735 -5920
rect -701 -5954 -638 -5920
rect -604 -5954 -539 -5920
rect -505 -5954 -442 -5920
rect -408 -5954 -343 -5920
rect -309 -5954 -246 -5920
rect -212 -5954 -147 -5920
rect -113 -5954 -50 -5920
rect -16 -5954 49 -5920
rect 83 -5954 146 -5920
rect 180 -5954 245 -5920
rect 279 -5954 342 -5920
rect 376 -5954 441 -5920
rect 475 -5954 538 -5920
rect 572 -5954 637 -5920
rect 671 -5954 734 -5920
rect 768 -5954 833 -5920
rect 867 -5954 930 -5920
rect 964 -5954 1029 -5920
rect 1063 -5954 1126 -5920
rect 1160 -5954 1225 -5920
rect 1259 -5954 1275 -5920
rect -1144 -5970 1275 -5954
rect -1130 -5992 -1090 -5970
rect -1032 -5992 -992 -5970
rect -934 -5992 -894 -5970
rect -836 -5992 -796 -5970
rect -738 -5992 -698 -5970
rect -640 -5992 -600 -5970
rect -542 -5992 -502 -5970
rect -444 -5992 -404 -5970
rect -346 -5992 -306 -5970
rect -248 -5992 -208 -5970
rect -150 -5992 -110 -5970
rect -52 -5992 -12 -5970
rect 46 -5992 86 -5970
rect 144 -5992 184 -5970
rect 242 -5992 282 -5970
rect 340 -5992 380 -5970
rect 438 -5992 478 -5970
rect 536 -5992 576 -5970
rect 634 -5992 674 -5970
rect 732 -5992 772 -5970
rect 830 -5992 870 -5970
rect 928 -5992 968 -5970
rect 1026 -5992 1066 -5970
rect 1124 -5992 1164 -5970
rect 1222 -5992 1262 -5970
rect -1130 -6414 -1090 -6392
rect -1032 -6414 -992 -6392
rect -934 -6414 -894 -6392
rect -836 -6414 -796 -6392
rect -738 -6414 -698 -6392
rect -640 -6414 -600 -6392
rect -542 -6414 -502 -6392
rect -444 -6414 -404 -6392
rect -346 -6414 -306 -6392
rect -248 -6414 -208 -6392
rect -150 -6414 -110 -6392
rect -52 -6414 -12 -6392
rect 46 -6414 86 -6392
rect 144 -6414 184 -6392
rect 242 -6414 282 -6392
rect 340 -6414 380 -6392
rect 438 -6414 478 -6392
rect 536 -6414 576 -6392
rect 634 -6414 674 -6392
rect 732 -6414 772 -6392
rect 830 -6414 870 -6392
rect 928 -6414 968 -6392
rect 1026 -6414 1066 -6392
rect 1124 -6414 1164 -6392
rect 1222 -6414 1262 -6392
rect -1144 -6430 1274 -6414
rect -1144 -6464 -1128 -6430
rect -1094 -6464 -1029 -6430
rect -995 -6464 -932 -6430
rect -898 -6464 -833 -6430
rect -799 -6464 -736 -6430
rect -702 -6464 -637 -6430
rect -603 -6464 -540 -6430
rect -506 -6464 -441 -6430
rect -407 -6464 -344 -6430
rect -310 -6464 -245 -6430
rect -211 -6464 -148 -6430
rect -114 -6464 -49 -6430
rect -15 -6464 48 -6430
rect 82 -6464 147 -6430
rect 181 -6464 244 -6430
rect 278 -6464 343 -6430
rect 377 -6464 440 -6430
rect 474 -6464 539 -6430
rect 573 -6464 636 -6430
rect 670 -6464 735 -6430
rect 769 -6464 832 -6430
rect 866 -6464 931 -6430
rect 965 -6464 1028 -6430
rect 1062 -6464 1127 -6430
rect 1161 -6464 1224 -6430
rect 1258 -6464 1274 -6430
rect -1144 -6480 1274 -6464
rect -1143 -6538 1275 -6522
rect -1143 -6572 -1127 -6538
rect -1093 -6572 -1029 -6538
rect -995 -6572 -931 -6538
rect -897 -6572 -833 -6538
rect -799 -6572 -735 -6538
rect -701 -6572 -637 -6538
rect -603 -6572 -539 -6538
rect -505 -6572 -441 -6538
rect -407 -6572 -343 -6538
rect -309 -6572 -245 -6538
rect -211 -6572 -147 -6538
rect -113 -6572 -49 -6538
rect -15 -6572 49 -6538
rect 83 -6572 147 -6538
rect 181 -6572 245 -6538
rect 279 -6572 343 -6538
rect 377 -6572 441 -6538
rect 475 -6572 539 -6538
rect 573 -6572 637 -6538
rect 671 -6572 735 -6538
rect 769 -6572 833 -6538
rect 867 -6572 931 -6538
rect 965 -6572 1029 -6538
rect 1063 -6572 1127 -6538
rect 1161 -6572 1225 -6538
rect 1259 -6572 1275 -6538
rect -1143 -6588 1275 -6572
rect -1130 -6610 -1090 -6588
rect -1032 -6610 -992 -6588
rect -934 -6610 -894 -6588
rect -836 -6610 -796 -6588
rect -738 -6610 -698 -6588
rect -640 -6610 -600 -6588
rect -542 -6610 -502 -6588
rect -444 -6610 -404 -6588
rect -346 -6610 -306 -6588
rect -248 -6610 -208 -6588
rect -150 -6610 -110 -6588
rect -52 -6610 -12 -6588
rect 46 -6610 86 -6588
rect 144 -6610 184 -6588
rect 242 -6610 282 -6588
rect 340 -6610 380 -6588
rect 438 -6610 478 -6588
rect 536 -6610 576 -6588
rect 634 -6610 674 -6588
rect 732 -6610 772 -6588
rect 830 -6610 870 -6588
rect 928 -6610 968 -6588
rect 1026 -6610 1066 -6588
rect 1124 -6610 1164 -6588
rect 1222 -6610 1262 -6588
rect -1130 -7032 -1090 -7010
rect -1032 -7032 -992 -7010
rect -934 -7032 -894 -7010
rect -836 -7032 -796 -7010
rect -738 -7032 -698 -7010
rect -640 -7032 -600 -7010
rect -542 -7032 -502 -7010
rect -444 -7032 -404 -7010
rect -346 -7032 -306 -7010
rect -248 -7032 -208 -7010
rect -150 -7032 -110 -7010
rect -52 -7032 -12 -7010
rect 46 -7032 86 -7010
rect 144 -7032 184 -7010
rect 242 -7032 282 -7010
rect 340 -7032 380 -7010
rect 438 -7032 478 -7010
rect 536 -7032 576 -7010
rect 634 -7032 674 -7010
rect 732 -7032 772 -7010
rect 830 -7032 870 -7010
rect 928 -7032 968 -7010
rect 1026 -7032 1066 -7010
rect 1124 -7032 1164 -7010
rect 1222 -7032 1262 -7010
rect -1143 -7048 1275 -7032
rect -1143 -7082 -1127 -7048
rect -1093 -7082 -1029 -7048
rect -995 -7082 -931 -7048
rect -897 -7082 -833 -7048
rect -799 -7082 -735 -7048
rect -701 -7082 -637 -7048
rect -603 -7082 -539 -7048
rect -505 -7082 -441 -7048
rect -407 -7082 -343 -7048
rect -309 -7082 -245 -7048
rect -211 -7082 -147 -7048
rect -113 -7082 -49 -7048
rect -15 -7082 49 -7048
rect 83 -7082 147 -7048
rect 181 -7082 245 -7048
rect 279 -7082 343 -7048
rect 377 -7082 441 -7048
rect 475 -7082 539 -7048
rect 573 -7082 637 -7048
rect 671 -7082 735 -7048
rect 769 -7082 833 -7048
rect 867 -7082 931 -7048
rect 965 -7082 1029 -7048
rect 1063 -7082 1127 -7048
rect 1161 -7082 1225 -7048
rect 1259 -7082 1275 -7048
rect -1143 -7098 1275 -7082
rect -1144 -7364 1275 -7348
rect -1144 -7398 -1127 -7364
rect -1093 -7398 -1030 -7364
rect -996 -7398 -931 -7364
rect -897 -7398 -834 -7364
rect -800 -7398 -735 -7364
rect -701 -7398 -638 -7364
rect -604 -7398 -539 -7364
rect -505 -7398 -442 -7364
rect -408 -7398 -343 -7364
rect -309 -7398 -246 -7364
rect -212 -7398 -147 -7364
rect -113 -7398 -50 -7364
rect -16 -7398 49 -7364
rect 83 -7398 146 -7364
rect 180 -7398 245 -7364
rect 279 -7398 342 -7364
rect 376 -7398 441 -7364
rect 475 -7398 538 -7364
rect 572 -7398 637 -7364
rect 671 -7398 734 -7364
rect 768 -7398 833 -7364
rect 867 -7398 930 -7364
rect 964 -7398 1029 -7364
rect 1063 -7398 1126 -7364
rect 1160 -7398 1225 -7364
rect 1259 -7398 1275 -7364
rect -1144 -7414 1275 -7398
rect -1130 -7436 -1090 -7414
rect -1032 -7436 -992 -7414
rect -934 -7436 -894 -7414
rect -836 -7436 -796 -7414
rect -738 -7436 -698 -7414
rect -640 -7436 -600 -7414
rect -542 -7436 -502 -7414
rect -444 -7436 -404 -7414
rect -346 -7436 -306 -7414
rect -248 -7436 -208 -7414
rect -150 -7436 -110 -7414
rect -52 -7436 -12 -7414
rect 46 -7436 86 -7414
rect 144 -7436 184 -7414
rect 242 -7436 282 -7414
rect 340 -7436 380 -7414
rect 438 -7436 478 -7414
rect 536 -7436 576 -7414
rect 634 -7436 674 -7414
rect 732 -7436 772 -7414
rect 830 -7436 870 -7414
rect 928 -7436 968 -7414
rect 1026 -7436 1066 -7414
rect 1124 -7436 1164 -7414
rect 1222 -7436 1262 -7414
rect -1130 -7858 -1090 -7836
rect -1032 -7858 -992 -7836
rect -934 -7858 -894 -7836
rect -836 -7858 -796 -7836
rect -738 -7858 -698 -7836
rect -640 -7858 -600 -7836
rect -542 -7858 -502 -7836
rect -444 -7858 -404 -7836
rect -346 -7858 -306 -7836
rect -248 -7858 -208 -7836
rect -150 -7858 -110 -7836
rect -52 -7858 -12 -7836
rect 46 -7858 86 -7836
rect 144 -7858 184 -7836
rect 242 -7858 282 -7836
rect 340 -7858 380 -7836
rect 438 -7858 478 -7836
rect 536 -7858 576 -7836
rect 634 -7858 674 -7836
rect 732 -7858 772 -7836
rect 830 -7858 870 -7836
rect 928 -7858 968 -7836
rect 1026 -7858 1066 -7836
rect 1124 -7858 1164 -7836
rect 1222 -7858 1262 -7836
rect -1144 -7874 1274 -7858
rect -1144 -7908 -1128 -7874
rect -1094 -7908 -1029 -7874
rect -995 -7908 -932 -7874
rect -898 -7908 -833 -7874
rect -799 -7908 -736 -7874
rect -702 -7908 -637 -7874
rect -603 -7908 -540 -7874
rect -506 -7908 -441 -7874
rect -407 -7908 -344 -7874
rect -310 -7908 -245 -7874
rect -211 -7908 -148 -7874
rect -114 -7908 -49 -7874
rect -15 -7908 48 -7874
rect 82 -7908 147 -7874
rect 181 -7908 244 -7874
rect 278 -7908 343 -7874
rect 377 -7908 440 -7874
rect 474 -7908 539 -7874
rect 573 -7908 636 -7874
rect 670 -7908 735 -7874
rect 769 -7908 832 -7874
rect 866 -7908 931 -7874
rect 965 -7908 1028 -7874
rect 1062 -7908 1127 -7874
rect 1161 -7908 1224 -7874
rect 1258 -7908 1274 -7874
rect -1144 -7924 1274 -7908
rect -1143 -7982 1275 -7966
rect -1143 -8016 -1127 -7982
rect -1093 -8016 -1029 -7982
rect -995 -8016 -931 -7982
rect -897 -8016 -833 -7982
rect -799 -8016 -735 -7982
rect -701 -8016 -637 -7982
rect -603 -8016 -539 -7982
rect -505 -8016 -441 -7982
rect -407 -8016 -343 -7982
rect -309 -8016 -245 -7982
rect -211 -8016 -147 -7982
rect -113 -8016 -49 -7982
rect -15 -8016 49 -7982
rect 83 -8016 147 -7982
rect 181 -8016 245 -7982
rect 279 -8016 343 -7982
rect 377 -8016 441 -7982
rect 475 -8016 539 -7982
rect 573 -8016 637 -7982
rect 671 -8016 735 -7982
rect 769 -8016 833 -7982
rect 867 -8016 931 -7982
rect 965 -8016 1029 -7982
rect 1063 -8016 1127 -7982
rect 1161 -8016 1225 -7982
rect 1259 -8016 1275 -7982
rect -1143 -8032 1275 -8016
rect -1130 -8054 -1090 -8032
rect -1032 -8054 -992 -8032
rect -934 -8054 -894 -8032
rect -836 -8054 -796 -8032
rect -738 -8054 -698 -8032
rect -640 -8054 -600 -8032
rect -542 -8054 -502 -8032
rect -444 -8054 -404 -8032
rect -346 -8054 -306 -8032
rect -248 -8054 -208 -8032
rect -150 -8054 -110 -8032
rect -52 -8054 -12 -8032
rect 46 -8054 86 -8032
rect 144 -8054 184 -8032
rect 242 -8054 282 -8032
rect 340 -8054 380 -8032
rect 438 -8054 478 -8032
rect 536 -8054 576 -8032
rect 634 -8054 674 -8032
rect 732 -8054 772 -8032
rect 830 -8054 870 -8032
rect 928 -8054 968 -8032
rect 1026 -8054 1066 -8032
rect 1124 -8054 1164 -8032
rect 1222 -8054 1262 -8032
rect -1130 -8476 -1090 -8454
rect -1032 -8476 -992 -8454
rect -934 -8476 -894 -8454
rect -836 -8476 -796 -8454
rect -738 -8476 -698 -8454
rect -640 -8476 -600 -8454
rect -542 -8476 -502 -8454
rect -444 -8476 -404 -8454
rect -346 -8476 -306 -8454
rect -248 -8476 -208 -8454
rect -150 -8476 -110 -8454
rect -52 -8476 -12 -8454
rect 46 -8476 86 -8454
rect 144 -8476 184 -8454
rect 242 -8476 282 -8454
rect 340 -8476 380 -8454
rect 438 -8476 478 -8454
rect 536 -8476 576 -8454
rect 634 -8476 674 -8454
rect 732 -8476 772 -8454
rect 830 -8476 870 -8454
rect 928 -8476 968 -8454
rect 1026 -8476 1066 -8454
rect 1124 -8476 1164 -8454
rect 1222 -8476 1262 -8454
rect -1143 -8492 1275 -8476
rect -1143 -8526 -1127 -8492
rect -1093 -8526 -1029 -8492
rect -995 -8526 -931 -8492
rect -897 -8526 -833 -8492
rect -799 -8526 -735 -8492
rect -701 -8526 -637 -8492
rect -603 -8526 -539 -8492
rect -505 -8526 -441 -8492
rect -407 -8526 -343 -8492
rect -309 -8526 -245 -8492
rect -211 -8526 -147 -8492
rect -113 -8526 -49 -8492
rect -15 -8526 49 -8492
rect 83 -8526 147 -8492
rect 181 -8526 245 -8492
rect 279 -8526 343 -8492
rect 377 -8526 441 -8492
rect 475 -8526 539 -8492
rect 573 -8526 637 -8492
rect 671 -8526 735 -8492
rect 769 -8526 833 -8492
rect 867 -8526 931 -8492
rect 965 -8526 1029 -8492
rect 1063 -8526 1127 -8492
rect 1161 -8526 1225 -8492
rect 1259 -8526 1275 -8492
rect -1143 -8542 1275 -8526
rect 2517 -6240 3955 -6224
rect 2517 -6274 2533 -6240
rect 2567 -6274 2631 -6240
rect 2665 -6274 2729 -6240
rect 2763 -6274 2827 -6240
rect 2861 -6274 2925 -6240
rect 2959 -6274 3023 -6240
rect 3057 -6274 3121 -6240
rect 3155 -6274 3219 -6240
rect 3253 -6274 3317 -6240
rect 3351 -6274 3415 -6240
rect 3449 -6274 3513 -6240
rect 3547 -6274 3611 -6240
rect 3645 -6274 3709 -6240
rect 3743 -6274 3807 -6240
rect 3841 -6274 3905 -6240
rect 3939 -6274 3955 -6240
rect 2517 -6290 3955 -6274
rect 2530 -6312 2570 -6290
rect 2628 -6312 2668 -6290
rect 2726 -6312 2766 -6290
rect 2824 -6312 2864 -6290
rect 2922 -6312 2962 -6290
rect 3020 -6312 3060 -6290
rect 3118 -6312 3158 -6290
rect 3216 -6312 3256 -6290
rect 3314 -6312 3354 -6290
rect 3412 -6312 3452 -6290
rect 3510 -6312 3550 -6290
rect 3608 -6312 3648 -6290
rect 3706 -6312 3746 -6290
rect 3804 -6312 3844 -6290
rect 3902 -6312 3942 -6290
rect 2530 -6734 2570 -6712
rect 2628 -6734 2668 -6712
rect 2726 -6734 2766 -6712
rect 2824 -6734 2864 -6712
rect 2922 -6734 2962 -6712
rect 3020 -6734 3060 -6712
rect 3118 -6734 3158 -6712
rect 3216 -6734 3256 -6712
rect 3314 -6734 3354 -6712
rect 3412 -6734 3452 -6712
rect 3510 -6734 3550 -6712
rect 3608 -6734 3648 -6712
rect 3706 -6734 3746 -6712
rect 3804 -6734 3844 -6712
rect 3902 -6734 3942 -6712
rect 2517 -6750 3955 -6734
rect 2517 -6784 2533 -6750
rect 2567 -6784 2631 -6750
rect 2665 -6784 2729 -6750
rect 2763 -6784 2827 -6750
rect 2861 -6784 2925 -6750
rect 2959 -6784 3023 -6750
rect 3057 -6784 3121 -6750
rect 3155 -6784 3219 -6750
rect 3253 -6784 3317 -6750
rect 3351 -6784 3415 -6750
rect 3449 -6784 3513 -6750
rect 3547 -6784 3611 -6750
rect 3645 -6784 3709 -6750
rect 3743 -6784 3807 -6750
rect 3841 -6784 3905 -6750
rect 3939 -6784 3955 -6750
rect 2517 -6800 3955 -6784
rect 2517 -6858 3955 -6842
rect 2517 -6892 2533 -6858
rect 2567 -6892 2631 -6858
rect 2665 -6892 2729 -6858
rect 2763 -6892 2827 -6858
rect 2861 -6892 2925 -6858
rect 2959 -6892 3023 -6858
rect 3057 -6892 3121 -6858
rect 3155 -6892 3219 -6858
rect 3253 -6892 3317 -6858
rect 3351 -6892 3415 -6858
rect 3449 -6892 3513 -6858
rect 3547 -6892 3611 -6858
rect 3645 -6892 3709 -6858
rect 3743 -6892 3807 -6858
rect 3841 -6892 3905 -6858
rect 3939 -6892 3955 -6858
rect 2517 -6908 3955 -6892
rect 2530 -6930 2570 -6908
rect 2628 -6930 2668 -6908
rect 2726 -6930 2766 -6908
rect 2824 -6930 2864 -6908
rect 2922 -6930 2962 -6908
rect 3020 -6930 3060 -6908
rect 3118 -6930 3158 -6908
rect 3216 -6930 3256 -6908
rect 3314 -6930 3354 -6908
rect 3412 -6930 3452 -6908
rect 3510 -6930 3550 -6908
rect 3608 -6930 3648 -6908
rect 3706 -6930 3746 -6908
rect 3804 -6930 3844 -6908
rect 3902 -6930 3942 -6908
rect 2530 -7352 2570 -7330
rect 2628 -7352 2668 -7330
rect 2726 -7352 2766 -7330
rect 2824 -7352 2864 -7330
rect 2922 -7352 2962 -7330
rect 3020 -7352 3060 -7330
rect 3118 -7352 3158 -7330
rect 3216 -7352 3256 -7330
rect 3314 -7352 3354 -7330
rect 3412 -7352 3452 -7330
rect 3510 -7352 3550 -7330
rect 3608 -7352 3648 -7330
rect 3706 -7352 3746 -7330
rect 3804 -7352 3844 -7330
rect 3902 -7352 3942 -7330
rect 2517 -7368 3955 -7352
rect 2517 -7402 2533 -7368
rect 2567 -7402 2631 -7368
rect 2665 -7402 2729 -7368
rect 2763 -7402 2827 -7368
rect 2861 -7402 2925 -7368
rect 2959 -7402 3023 -7368
rect 3057 -7402 3121 -7368
rect 3155 -7402 3219 -7368
rect 3253 -7402 3317 -7368
rect 3351 -7402 3415 -7368
rect 3449 -7402 3513 -7368
rect 3547 -7402 3611 -7368
rect 3645 -7402 3709 -7368
rect 3743 -7402 3807 -7368
rect 3841 -7402 3905 -7368
rect 3939 -7402 3955 -7368
rect 2517 -7418 3955 -7402
rect 1646 -8018 2768 -8002
rect 1646 -8052 1662 -8018
rect 1696 -8052 1758 -8018
rect 1792 -8052 1854 -8018
rect 1888 -8052 1950 -8018
rect 1984 -8052 2046 -8018
rect 2080 -8052 2142 -8018
rect 2176 -8052 2238 -8018
rect 2272 -8052 2334 -8018
rect 2368 -8052 2430 -8018
rect 2464 -8052 2526 -8018
rect 2560 -8052 2622 -8018
rect 2656 -8052 2718 -8018
rect 2752 -8052 2768 -8018
rect 1646 -8068 2768 -8052
rect 1664 -8090 1694 -8068
rect 1760 -8090 1790 -8068
rect 1856 -8090 1886 -8068
rect 1952 -8090 1982 -8068
rect 2048 -8090 2078 -8068
rect 2144 -8090 2174 -8068
rect 2240 -8090 2270 -8068
rect 2336 -8090 2366 -8068
rect 2432 -8090 2462 -8068
rect 2528 -8090 2558 -8068
rect 2624 -8090 2654 -8068
rect 2720 -8090 2750 -8068
rect 1664 -8512 1694 -8490
rect 1760 -8512 1790 -8490
rect 1856 -8512 1886 -8490
rect 1952 -8512 1982 -8490
rect 2048 -8512 2078 -8490
rect 2144 -8512 2174 -8490
rect 2240 -8512 2270 -8490
rect 2336 -8512 2366 -8490
rect 2432 -8512 2462 -8490
rect 2528 -8512 2558 -8490
rect 2624 -8512 2654 -8490
rect 2720 -8512 2750 -8490
rect 1646 -8528 2768 -8512
rect 1646 -8562 1662 -8528
rect 1696 -8562 1758 -8528
rect 1792 -8562 1854 -8528
rect 1888 -8562 1950 -8528
rect 1984 -8562 2046 -8528
rect 2080 -8562 2142 -8528
rect 2176 -8562 2238 -8528
rect 2272 -8562 2334 -8528
rect 2368 -8562 2430 -8528
rect 2464 -8562 2526 -8528
rect 2560 -8562 2622 -8528
rect 2656 -8562 2718 -8528
rect 2752 -8562 2768 -8528
rect 1646 -8578 2768 -8562
rect 3542 -8018 4664 -8002
rect 3542 -8052 3558 -8018
rect 3592 -8052 3654 -8018
rect 3688 -8052 3750 -8018
rect 3784 -8052 3846 -8018
rect 3880 -8052 3942 -8018
rect 3976 -8052 4038 -8018
rect 4072 -8052 4134 -8018
rect 4168 -8052 4230 -8018
rect 4264 -8052 4326 -8018
rect 4360 -8052 4422 -8018
rect 4456 -8052 4518 -8018
rect 4552 -8052 4614 -8018
rect 4648 -8052 4664 -8018
rect 3542 -8068 4664 -8052
rect 3560 -8090 3590 -8068
rect 3656 -8090 3686 -8068
rect 3752 -8090 3782 -8068
rect 3848 -8090 3878 -8068
rect 3944 -8090 3974 -8068
rect 4040 -8090 4070 -8068
rect 4136 -8090 4166 -8068
rect 4232 -8090 4262 -8068
rect 4328 -8090 4358 -8068
rect 4424 -8090 4454 -8068
rect 4520 -8090 4550 -8068
rect 4616 -8090 4646 -8068
rect 3560 -8512 3590 -8490
rect 3656 -8512 3686 -8490
rect 3752 -8512 3782 -8490
rect 3848 -8512 3878 -8490
rect 3944 -8512 3974 -8490
rect 4040 -8512 4070 -8490
rect 4136 -8512 4166 -8490
rect 4232 -8512 4262 -8490
rect 4328 -8512 4358 -8490
rect 4424 -8512 4454 -8490
rect 4520 -8512 4550 -8490
rect 4616 -8512 4646 -8490
rect 3542 -8528 4664 -8512
rect 3542 -8562 3558 -8528
rect 3592 -8562 3654 -8528
rect 3688 -8562 3750 -8528
rect 3784 -8562 3846 -8528
rect 3880 -8562 3942 -8528
rect 3976 -8562 4038 -8528
rect 4072 -8562 4134 -8528
rect 4168 -8562 4230 -8528
rect 4264 -8562 4326 -8528
rect 4360 -8562 4422 -8528
rect 4456 -8562 4518 -8528
rect 4552 -8562 4614 -8528
rect 4648 -8562 4664 -8528
rect 3542 -8578 4664 -8562
rect -1164 -8784 -1098 -8768
rect -1164 -8818 -1148 -8784
rect -1114 -8818 -1098 -8784
rect -1164 -8834 -1098 -8818
rect -972 -8784 -906 -8768
rect -972 -8818 -956 -8784
rect -922 -8818 -906 -8784
rect -1146 -8856 -1116 -8834
rect -1050 -8856 -1020 -8830
rect -972 -8834 -906 -8818
rect -780 -8784 -714 -8768
rect -780 -8818 -764 -8784
rect -730 -8818 -714 -8784
rect -954 -8856 -924 -8834
rect -858 -8856 -828 -8830
rect -780 -8834 -714 -8818
rect -588 -8784 -522 -8768
rect -588 -8818 -572 -8784
rect -538 -8818 -522 -8784
rect -762 -8856 -732 -8834
rect -666 -8856 -636 -8830
rect -588 -8834 -522 -8818
rect -396 -8784 -330 -8768
rect -396 -8818 -380 -8784
rect -346 -8818 -330 -8784
rect -570 -8856 -540 -8834
rect -474 -8856 -444 -8830
rect -396 -8834 -330 -8818
rect -204 -8784 -138 -8768
rect -204 -8818 -188 -8784
rect -154 -8818 -138 -8784
rect -378 -8856 -348 -8834
rect -282 -8856 -252 -8830
rect -204 -8834 -138 -8818
rect -12 -8784 54 -8768
rect -12 -8818 4 -8784
rect 38 -8818 54 -8784
rect -186 -8856 -156 -8834
rect -90 -8856 -60 -8830
rect -12 -8834 54 -8818
rect 180 -8784 246 -8768
rect 180 -8818 196 -8784
rect 230 -8818 246 -8784
rect 6 -8856 36 -8834
rect 102 -8856 132 -8830
rect 180 -8834 246 -8818
rect 372 -8784 438 -8768
rect 372 -8818 388 -8784
rect 422 -8818 438 -8784
rect 198 -8856 228 -8834
rect 294 -8856 324 -8830
rect 372 -8834 438 -8818
rect 564 -8784 630 -8768
rect 564 -8818 580 -8784
rect 614 -8818 630 -8784
rect 390 -8856 420 -8834
rect 486 -8856 516 -8830
rect 564 -8834 630 -8818
rect 756 -8784 822 -8768
rect 756 -8818 772 -8784
rect 806 -8818 822 -8784
rect 582 -8856 612 -8834
rect 678 -8856 708 -8830
rect 756 -8834 822 -8818
rect 948 -8784 1014 -8768
rect 948 -8818 964 -8784
rect 998 -8818 1014 -8784
rect 774 -8856 804 -8834
rect 870 -8856 900 -8830
rect 948 -8834 1014 -8818
rect 1140 -8784 1206 -8768
rect 1140 -8818 1156 -8784
rect 1190 -8818 1206 -8784
rect 966 -8856 996 -8834
rect 1062 -8856 1092 -8830
rect 1140 -8834 1206 -8818
rect 1158 -8856 1188 -8834
rect -1146 -9282 -1116 -9256
rect -1050 -9278 -1020 -9256
rect -1068 -9294 -1002 -9278
rect -954 -9282 -924 -9256
rect -858 -9278 -828 -9256
rect -1068 -9328 -1052 -9294
rect -1018 -9328 -1002 -9294
rect -1068 -9344 -1002 -9328
rect -876 -9294 -810 -9278
rect -762 -9282 -732 -9256
rect -666 -9278 -636 -9256
rect -876 -9328 -860 -9294
rect -826 -9328 -810 -9294
rect -876 -9344 -810 -9328
rect -684 -9294 -618 -9278
rect -570 -9282 -540 -9256
rect -474 -9278 -444 -9256
rect -684 -9328 -668 -9294
rect -634 -9328 -618 -9294
rect -684 -9344 -618 -9328
rect -492 -9294 -426 -9278
rect -378 -9282 -348 -9256
rect -282 -9278 -252 -9256
rect -492 -9328 -476 -9294
rect -442 -9328 -426 -9294
rect -492 -9344 -426 -9328
rect -300 -9294 -234 -9278
rect -186 -9282 -156 -9256
rect -90 -9278 -60 -9256
rect -300 -9328 -284 -9294
rect -250 -9328 -234 -9294
rect -300 -9344 -234 -9328
rect -108 -9294 -42 -9278
rect 6 -9282 36 -9256
rect 102 -9278 132 -9256
rect -108 -9328 -92 -9294
rect -58 -9328 -42 -9294
rect -108 -9344 -42 -9328
rect 84 -9294 150 -9278
rect 198 -9282 228 -9256
rect 294 -9278 324 -9256
rect 84 -9328 100 -9294
rect 134 -9328 150 -9294
rect 84 -9344 150 -9328
rect 276 -9294 342 -9278
rect 390 -9282 420 -9256
rect 486 -9278 516 -9256
rect 276 -9328 292 -9294
rect 326 -9328 342 -9294
rect 276 -9344 342 -9328
rect 468 -9294 534 -9278
rect 582 -9282 612 -9256
rect 678 -9278 708 -9256
rect 468 -9328 484 -9294
rect 518 -9328 534 -9294
rect 468 -9344 534 -9328
rect 660 -9294 726 -9278
rect 774 -9282 804 -9256
rect 870 -9278 900 -9256
rect 660 -9328 676 -9294
rect 710 -9328 726 -9294
rect 660 -9344 726 -9328
rect 852 -9294 918 -9278
rect 966 -9282 996 -9256
rect 1062 -9278 1092 -9256
rect 852 -9328 868 -9294
rect 902 -9328 918 -9294
rect 852 -9344 918 -9328
rect 1044 -9294 1110 -9278
rect 1158 -9282 1188 -9256
rect 1044 -9328 1060 -9294
rect 1094 -9328 1110 -9294
rect 1044 -9344 1110 -9328
rect -1068 -9402 -1002 -9386
rect -1068 -9436 -1052 -9402
rect -1018 -9436 -1002 -9402
rect -1146 -9474 -1116 -9448
rect -1068 -9452 -1002 -9436
rect -876 -9402 -810 -9386
rect -876 -9436 -860 -9402
rect -826 -9436 -810 -9402
rect -1050 -9474 -1020 -9452
rect -954 -9474 -924 -9448
rect -876 -9452 -810 -9436
rect -684 -9402 -618 -9386
rect -684 -9436 -668 -9402
rect -634 -9436 -618 -9402
rect -858 -9474 -828 -9452
rect -762 -9474 -732 -9448
rect -684 -9452 -618 -9436
rect -492 -9402 -426 -9386
rect -492 -9436 -476 -9402
rect -442 -9436 -426 -9402
rect -666 -9474 -636 -9452
rect -570 -9474 -540 -9448
rect -492 -9452 -426 -9436
rect -300 -9402 -234 -9386
rect -300 -9436 -284 -9402
rect -250 -9436 -234 -9402
rect -474 -9474 -444 -9452
rect -378 -9474 -348 -9448
rect -300 -9452 -234 -9436
rect -108 -9402 -42 -9386
rect -108 -9436 -92 -9402
rect -58 -9436 -42 -9402
rect -282 -9474 -252 -9452
rect -186 -9474 -156 -9448
rect -108 -9452 -42 -9436
rect 84 -9402 150 -9386
rect 84 -9436 100 -9402
rect 134 -9436 150 -9402
rect -90 -9474 -60 -9452
rect 6 -9474 36 -9448
rect 84 -9452 150 -9436
rect 276 -9402 342 -9386
rect 276 -9436 292 -9402
rect 326 -9436 342 -9402
rect 102 -9474 132 -9452
rect 198 -9474 228 -9448
rect 276 -9452 342 -9436
rect 468 -9402 534 -9386
rect 468 -9436 484 -9402
rect 518 -9436 534 -9402
rect 294 -9474 324 -9452
rect 390 -9474 420 -9448
rect 468 -9452 534 -9436
rect 660 -9402 726 -9386
rect 660 -9436 676 -9402
rect 710 -9436 726 -9402
rect 486 -9474 516 -9452
rect 582 -9474 612 -9448
rect 660 -9452 726 -9436
rect 852 -9402 918 -9386
rect 852 -9436 868 -9402
rect 902 -9436 918 -9402
rect 678 -9474 708 -9452
rect 774 -9474 804 -9448
rect 852 -9452 918 -9436
rect 1044 -9402 1110 -9386
rect 1044 -9436 1060 -9402
rect 1094 -9436 1110 -9402
rect 870 -9474 900 -9452
rect 966 -9474 996 -9448
rect 1044 -9452 1110 -9436
rect 1062 -9474 1092 -9452
rect 1158 -9474 1188 -9448
rect -1146 -9896 -1116 -9874
rect -1164 -9912 -1098 -9896
rect -1050 -9900 -1020 -9874
rect -954 -9896 -924 -9874
rect -1164 -9946 -1148 -9912
rect -1114 -9946 -1098 -9912
rect -1164 -9962 -1098 -9946
rect -972 -9912 -906 -9896
rect -858 -9900 -828 -9874
rect -762 -9896 -732 -9874
rect -972 -9946 -956 -9912
rect -922 -9946 -906 -9912
rect -972 -9962 -906 -9946
rect -780 -9912 -714 -9896
rect -666 -9900 -636 -9874
rect -570 -9896 -540 -9874
rect -780 -9946 -764 -9912
rect -730 -9946 -714 -9912
rect -780 -9962 -714 -9946
rect -588 -9912 -522 -9896
rect -474 -9900 -444 -9874
rect -378 -9896 -348 -9874
rect -588 -9946 -572 -9912
rect -538 -9946 -522 -9912
rect -588 -9962 -522 -9946
rect -396 -9912 -330 -9896
rect -282 -9900 -252 -9874
rect -186 -9896 -156 -9874
rect -396 -9946 -380 -9912
rect -346 -9946 -330 -9912
rect -396 -9962 -330 -9946
rect -204 -9912 -138 -9896
rect -90 -9900 -60 -9874
rect 6 -9896 36 -9874
rect -204 -9946 -188 -9912
rect -154 -9946 -138 -9912
rect -204 -9962 -138 -9946
rect -12 -9912 54 -9896
rect 102 -9900 132 -9874
rect 198 -9896 228 -9874
rect -12 -9946 4 -9912
rect 38 -9946 54 -9912
rect -12 -9962 54 -9946
rect 180 -9912 246 -9896
rect 294 -9900 324 -9874
rect 390 -9896 420 -9874
rect 180 -9946 196 -9912
rect 230 -9946 246 -9912
rect 180 -9962 246 -9946
rect 372 -9912 438 -9896
rect 486 -9900 516 -9874
rect 582 -9896 612 -9874
rect 372 -9946 388 -9912
rect 422 -9946 438 -9912
rect 372 -9962 438 -9946
rect 564 -9912 630 -9896
rect 678 -9900 708 -9874
rect 774 -9896 804 -9874
rect 564 -9946 580 -9912
rect 614 -9946 630 -9912
rect 564 -9962 630 -9946
rect 756 -9912 822 -9896
rect 870 -9900 900 -9874
rect 966 -9896 996 -9874
rect 756 -9946 772 -9912
rect 806 -9946 822 -9912
rect 756 -9962 822 -9946
rect 948 -9912 1014 -9896
rect 1062 -9900 1092 -9874
rect 1158 -9896 1188 -9874
rect 948 -9946 964 -9912
rect 998 -9946 1014 -9912
rect 948 -9962 1014 -9946
rect 1140 -9912 1206 -9896
rect 1140 -9946 1156 -9912
rect 1190 -9946 1206 -9912
rect 1140 -9962 1206 -9946
rect -1164 -10020 -1098 -10004
rect -1164 -10054 -1148 -10020
rect -1114 -10054 -1098 -10020
rect -1164 -10070 -1098 -10054
rect -972 -10020 -906 -10004
rect -972 -10054 -956 -10020
rect -922 -10054 -906 -10020
rect -1146 -10092 -1116 -10070
rect -1050 -10092 -1020 -10066
rect -972 -10070 -906 -10054
rect -780 -10020 -714 -10004
rect -780 -10054 -764 -10020
rect -730 -10054 -714 -10020
rect -954 -10092 -924 -10070
rect -858 -10092 -828 -10066
rect -780 -10070 -714 -10054
rect -588 -10020 -522 -10004
rect -588 -10054 -572 -10020
rect -538 -10054 -522 -10020
rect -762 -10092 -732 -10070
rect -666 -10092 -636 -10066
rect -588 -10070 -522 -10054
rect -396 -10020 -330 -10004
rect -396 -10054 -380 -10020
rect -346 -10054 -330 -10020
rect -570 -10092 -540 -10070
rect -474 -10092 -444 -10066
rect -396 -10070 -330 -10054
rect -204 -10020 -138 -10004
rect -204 -10054 -188 -10020
rect -154 -10054 -138 -10020
rect -378 -10092 -348 -10070
rect -282 -10092 -252 -10066
rect -204 -10070 -138 -10054
rect -12 -10020 54 -10004
rect -12 -10054 4 -10020
rect 38 -10054 54 -10020
rect -186 -10092 -156 -10070
rect -90 -10092 -60 -10066
rect -12 -10070 54 -10054
rect 180 -10020 246 -10004
rect 180 -10054 196 -10020
rect 230 -10054 246 -10020
rect 6 -10092 36 -10070
rect 102 -10092 132 -10066
rect 180 -10070 246 -10054
rect 372 -10020 438 -10004
rect 372 -10054 388 -10020
rect 422 -10054 438 -10020
rect 198 -10092 228 -10070
rect 294 -10092 324 -10066
rect 372 -10070 438 -10054
rect 564 -10020 630 -10004
rect 564 -10054 580 -10020
rect 614 -10054 630 -10020
rect 390 -10092 420 -10070
rect 486 -10092 516 -10066
rect 564 -10070 630 -10054
rect 756 -10020 822 -10004
rect 756 -10054 772 -10020
rect 806 -10054 822 -10020
rect 582 -10092 612 -10070
rect 678 -10092 708 -10066
rect 756 -10070 822 -10054
rect 948 -10020 1014 -10004
rect 948 -10054 964 -10020
rect 998 -10054 1014 -10020
rect 774 -10092 804 -10070
rect 870 -10092 900 -10066
rect 948 -10070 1014 -10054
rect 1140 -10020 1206 -10004
rect 1140 -10054 1156 -10020
rect 1190 -10054 1206 -10020
rect 966 -10092 996 -10070
rect 1062 -10092 1092 -10066
rect 1140 -10070 1206 -10054
rect 1158 -10092 1188 -10070
rect -1146 -10518 -1116 -10492
rect -1050 -10514 -1020 -10492
rect -1068 -10530 -1002 -10514
rect -954 -10518 -924 -10492
rect -858 -10514 -828 -10492
rect -1068 -10564 -1052 -10530
rect -1018 -10564 -1002 -10530
rect -1068 -10580 -1002 -10564
rect -876 -10530 -810 -10514
rect -762 -10518 -732 -10492
rect -666 -10514 -636 -10492
rect -876 -10564 -860 -10530
rect -826 -10564 -810 -10530
rect -876 -10580 -810 -10564
rect -684 -10530 -618 -10514
rect -570 -10518 -540 -10492
rect -474 -10514 -444 -10492
rect -684 -10564 -668 -10530
rect -634 -10564 -618 -10530
rect -684 -10580 -618 -10564
rect -492 -10530 -426 -10514
rect -378 -10518 -348 -10492
rect -282 -10514 -252 -10492
rect -492 -10564 -476 -10530
rect -442 -10564 -426 -10530
rect -492 -10580 -426 -10564
rect -300 -10530 -234 -10514
rect -186 -10518 -156 -10492
rect -90 -10514 -60 -10492
rect -300 -10564 -284 -10530
rect -250 -10564 -234 -10530
rect -300 -10580 -234 -10564
rect -108 -10530 -42 -10514
rect 6 -10518 36 -10492
rect 102 -10514 132 -10492
rect -108 -10564 -92 -10530
rect -58 -10564 -42 -10530
rect -108 -10580 -42 -10564
rect 84 -10530 150 -10514
rect 198 -10518 228 -10492
rect 294 -10514 324 -10492
rect 84 -10564 100 -10530
rect 134 -10564 150 -10530
rect 84 -10580 150 -10564
rect 276 -10530 342 -10514
rect 390 -10518 420 -10492
rect 486 -10514 516 -10492
rect 276 -10564 292 -10530
rect 326 -10564 342 -10530
rect 276 -10580 342 -10564
rect 468 -10530 534 -10514
rect 582 -10518 612 -10492
rect 678 -10514 708 -10492
rect 468 -10564 484 -10530
rect 518 -10564 534 -10530
rect 468 -10580 534 -10564
rect 660 -10530 726 -10514
rect 774 -10518 804 -10492
rect 870 -10514 900 -10492
rect 660 -10564 676 -10530
rect 710 -10564 726 -10530
rect 660 -10580 726 -10564
rect 852 -10530 918 -10514
rect 966 -10518 996 -10492
rect 1062 -10514 1092 -10492
rect 852 -10564 868 -10530
rect 902 -10564 918 -10530
rect 852 -10580 918 -10564
rect 1044 -10530 1110 -10514
rect 1158 -10518 1188 -10492
rect 1044 -10564 1060 -10530
rect 1094 -10564 1110 -10530
rect 1044 -10580 1110 -10564
rect -1068 -10638 -1002 -10622
rect -1068 -10672 -1052 -10638
rect -1018 -10672 -1002 -10638
rect -1146 -10710 -1116 -10684
rect -1068 -10688 -1002 -10672
rect -876 -10638 -810 -10622
rect -876 -10672 -860 -10638
rect -826 -10672 -810 -10638
rect -1050 -10710 -1020 -10688
rect -954 -10710 -924 -10684
rect -876 -10688 -810 -10672
rect -684 -10638 -618 -10622
rect -684 -10672 -668 -10638
rect -634 -10672 -618 -10638
rect -858 -10710 -828 -10688
rect -762 -10710 -732 -10684
rect -684 -10688 -618 -10672
rect -492 -10638 -426 -10622
rect -492 -10672 -476 -10638
rect -442 -10672 -426 -10638
rect -666 -10710 -636 -10688
rect -570 -10710 -540 -10684
rect -492 -10688 -426 -10672
rect -300 -10638 -234 -10622
rect -300 -10672 -284 -10638
rect -250 -10672 -234 -10638
rect -474 -10710 -444 -10688
rect -378 -10710 -348 -10684
rect -300 -10688 -234 -10672
rect -108 -10638 -42 -10622
rect -108 -10672 -92 -10638
rect -58 -10672 -42 -10638
rect -282 -10710 -252 -10688
rect -186 -10710 -156 -10684
rect -108 -10688 -42 -10672
rect 84 -10638 150 -10622
rect 84 -10672 100 -10638
rect 134 -10672 150 -10638
rect -90 -10710 -60 -10688
rect 6 -10710 36 -10684
rect 84 -10688 150 -10672
rect 276 -10638 342 -10622
rect 276 -10672 292 -10638
rect 326 -10672 342 -10638
rect 102 -10710 132 -10688
rect 198 -10710 228 -10684
rect 276 -10688 342 -10672
rect 468 -10638 534 -10622
rect 468 -10672 484 -10638
rect 518 -10672 534 -10638
rect 294 -10710 324 -10688
rect 390 -10710 420 -10684
rect 468 -10688 534 -10672
rect 660 -10638 726 -10622
rect 660 -10672 676 -10638
rect 710 -10672 726 -10638
rect 486 -10710 516 -10688
rect 582 -10710 612 -10684
rect 660 -10688 726 -10672
rect 852 -10638 918 -10622
rect 852 -10672 868 -10638
rect 902 -10672 918 -10638
rect 678 -10710 708 -10688
rect 774 -10710 804 -10684
rect 852 -10688 918 -10672
rect 1044 -10638 1110 -10622
rect 1044 -10672 1060 -10638
rect 1094 -10672 1110 -10638
rect 870 -10710 900 -10688
rect 966 -10710 996 -10684
rect 1044 -10688 1110 -10672
rect 1062 -10710 1092 -10688
rect 1158 -10710 1188 -10684
rect -1146 -11132 -1116 -11110
rect -1164 -11148 -1098 -11132
rect -1050 -11136 -1020 -11110
rect -954 -11132 -924 -11110
rect -1164 -11182 -1148 -11148
rect -1114 -11182 -1098 -11148
rect -1164 -11198 -1098 -11182
rect -972 -11148 -906 -11132
rect -858 -11136 -828 -11110
rect -762 -11132 -732 -11110
rect -972 -11182 -956 -11148
rect -922 -11182 -906 -11148
rect -972 -11198 -906 -11182
rect -780 -11148 -714 -11132
rect -666 -11136 -636 -11110
rect -570 -11132 -540 -11110
rect -780 -11182 -764 -11148
rect -730 -11182 -714 -11148
rect -780 -11198 -714 -11182
rect -588 -11148 -522 -11132
rect -474 -11136 -444 -11110
rect -378 -11132 -348 -11110
rect -588 -11182 -572 -11148
rect -538 -11182 -522 -11148
rect -588 -11198 -522 -11182
rect -396 -11148 -330 -11132
rect -282 -11136 -252 -11110
rect -186 -11132 -156 -11110
rect -396 -11182 -380 -11148
rect -346 -11182 -330 -11148
rect -396 -11198 -330 -11182
rect -204 -11148 -138 -11132
rect -90 -11136 -60 -11110
rect 6 -11132 36 -11110
rect -204 -11182 -188 -11148
rect -154 -11182 -138 -11148
rect -204 -11198 -138 -11182
rect -12 -11148 54 -11132
rect 102 -11136 132 -11110
rect 198 -11132 228 -11110
rect -12 -11182 4 -11148
rect 38 -11182 54 -11148
rect -12 -11198 54 -11182
rect 180 -11148 246 -11132
rect 294 -11136 324 -11110
rect 390 -11132 420 -11110
rect 180 -11182 196 -11148
rect 230 -11182 246 -11148
rect 180 -11198 246 -11182
rect 372 -11148 438 -11132
rect 486 -11136 516 -11110
rect 582 -11132 612 -11110
rect 372 -11182 388 -11148
rect 422 -11182 438 -11148
rect 372 -11198 438 -11182
rect 564 -11148 630 -11132
rect 678 -11136 708 -11110
rect 774 -11132 804 -11110
rect 564 -11182 580 -11148
rect 614 -11182 630 -11148
rect 564 -11198 630 -11182
rect 756 -11148 822 -11132
rect 870 -11136 900 -11110
rect 966 -11132 996 -11110
rect 756 -11182 772 -11148
rect 806 -11182 822 -11148
rect 756 -11198 822 -11182
rect 948 -11148 1014 -11132
rect 1062 -11136 1092 -11110
rect 1158 -11132 1188 -11110
rect 948 -11182 964 -11148
rect 998 -11182 1014 -11148
rect 948 -11198 1014 -11182
rect 1140 -11148 1206 -11132
rect 1140 -11182 1156 -11148
rect 1190 -11182 1206 -11148
rect 1140 -11198 1206 -11182
rect 1660 -8838 1860 -8822
rect 1660 -8872 1676 -8838
rect 1844 -8872 1860 -8838
rect 1660 -8910 1860 -8872
rect 1918 -8838 2118 -8822
rect 1918 -8872 1934 -8838
rect 2102 -8872 2118 -8838
rect 1918 -8910 2118 -8872
rect 2176 -8838 2376 -8822
rect 2176 -8872 2192 -8838
rect 2360 -8872 2376 -8838
rect 2176 -8910 2376 -8872
rect 2434 -8838 2634 -8822
rect 2434 -8872 2450 -8838
rect 2618 -8872 2634 -8838
rect 2434 -8910 2634 -8872
rect 2692 -8838 2892 -8822
rect 2692 -8872 2708 -8838
rect 2876 -8872 2892 -8838
rect 2692 -8910 2892 -8872
rect 2950 -8838 3150 -8822
rect 2950 -8872 2966 -8838
rect 3134 -8872 3150 -8838
rect 2950 -8910 3150 -8872
rect 1660 -9348 1860 -9310
rect 1660 -9382 1676 -9348
rect 1844 -9382 1860 -9348
rect 1660 -9398 1860 -9382
rect 1918 -9348 2118 -9310
rect 1918 -9382 1934 -9348
rect 2102 -9382 2118 -9348
rect 1918 -9398 2118 -9382
rect 2176 -9348 2376 -9310
rect 2176 -9382 2192 -9348
rect 2360 -9382 2376 -9348
rect 2176 -9398 2376 -9382
rect 2434 -9348 2634 -9310
rect 2434 -9382 2450 -9348
rect 2618 -9382 2634 -9348
rect 2434 -9398 2634 -9382
rect 2692 -9348 2892 -9310
rect 2692 -9382 2708 -9348
rect 2876 -9382 2892 -9348
rect 2692 -9398 2892 -9382
rect 2950 -9348 3150 -9310
rect 2950 -9382 2966 -9348
rect 3134 -9382 3150 -9348
rect 2950 -9398 3150 -9382
rect 3556 -8838 3756 -8822
rect 3556 -8872 3572 -8838
rect 3740 -8872 3756 -8838
rect 3556 -8910 3756 -8872
rect 3814 -8838 4014 -8822
rect 3814 -8872 3830 -8838
rect 3998 -8872 4014 -8838
rect 3814 -8910 4014 -8872
rect 4072 -8838 4272 -8822
rect 4072 -8872 4088 -8838
rect 4256 -8872 4272 -8838
rect 4072 -8910 4272 -8872
rect 4330 -8838 4530 -8822
rect 4330 -8872 4346 -8838
rect 4514 -8872 4530 -8838
rect 4330 -8910 4530 -8872
rect 4588 -8838 4788 -8822
rect 4588 -8872 4604 -8838
rect 4772 -8872 4788 -8838
rect 4588 -8910 4788 -8872
rect 4846 -8838 5046 -8822
rect 4846 -8872 4862 -8838
rect 5030 -8872 5046 -8838
rect 4846 -8910 5046 -8872
rect 3556 -9348 3756 -9310
rect 3556 -9382 3572 -9348
rect 3740 -9382 3756 -9348
rect 3556 -9398 3756 -9382
rect 3814 -9348 4014 -9310
rect 3814 -9382 3830 -9348
rect 3998 -9382 4014 -9348
rect 3814 -9398 4014 -9382
rect 4072 -9348 4272 -9310
rect 4072 -9382 4088 -9348
rect 4256 -9382 4272 -9348
rect 4072 -9398 4272 -9382
rect 4330 -9348 4530 -9310
rect 4330 -9382 4346 -9348
rect 4514 -9382 4530 -9348
rect 4330 -9398 4530 -9382
rect 4588 -9348 4788 -9310
rect 4588 -9382 4604 -9348
rect 4772 -9382 4788 -9348
rect 4588 -9398 4788 -9382
rect 4846 -9348 5046 -9310
rect 4846 -9382 4862 -9348
rect 5030 -9382 5046 -9348
rect 4846 -9398 5046 -9382
rect 5588 -8838 5654 -8822
rect 5588 -8872 5604 -8838
rect 5638 -8872 5654 -8838
rect 5510 -8910 5540 -8884
rect 5588 -8888 5654 -8872
rect 5780 -8838 5846 -8822
rect 5780 -8872 5796 -8838
rect 5830 -8872 5846 -8838
rect 5606 -8910 5636 -8888
rect 5702 -8910 5732 -8884
rect 5780 -8888 5846 -8872
rect 5798 -8910 5828 -8888
rect 5894 -8910 5924 -8884
rect 5510 -9332 5540 -9310
rect 5492 -9348 5558 -9332
rect 5606 -9336 5636 -9310
rect 5702 -9332 5732 -9310
rect 5492 -9382 5508 -9348
rect 5542 -9382 5558 -9348
rect 5492 -9398 5558 -9382
rect 5684 -9348 5750 -9332
rect 5798 -9336 5828 -9310
rect 5894 -9332 5924 -9310
rect 5684 -9382 5700 -9348
rect 5734 -9382 5750 -9348
rect 5684 -9398 5750 -9382
rect 5876 -9348 5942 -9332
rect 5876 -9382 5892 -9348
rect 5926 -9382 5942 -9348
rect 5876 -9398 5942 -9382
rect 1693 -9850 2093 -9834
rect 1693 -9884 1709 -9850
rect 2077 -9884 2093 -9850
rect 1693 -9922 2093 -9884
rect 2613 -9850 3013 -9834
rect 2613 -9884 2629 -9850
rect 2997 -9884 3013 -9850
rect 2613 -9922 3013 -9884
rect 3533 -9850 3933 -9834
rect 3533 -9884 3549 -9850
rect 3917 -9884 3933 -9850
rect 3533 -9922 3933 -9884
rect 4453 -9850 4853 -9834
rect 4453 -9884 4469 -9850
rect 4837 -9884 4853 -9850
rect 4453 -9922 4853 -9884
rect 5373 -9850 5773 -9834
rect 5373 -9884 5389 -9850
rect 5757 -9884 5773 -9850
rect 5373 -9922 5773 -9884
rect 1693 -10960 2093 -10922
rect 1693 -10994 1709 -10960
rect 2077 -10994 2093 -10960
rect 1693 -11010 2093 -10994
rect 2613 -10960 3013 -10922
rect 2613 -10994 2629 -10960
rect 2997 -10994 3013 -10960
rect 2613 -11010 3013 -10994
rect 3533 -10960 3933 -10922
rect 3533 -10994 3549 -10960
rect 3917 -10994 3933 -10960
rect 3533 -11010 3933 -10994
rect 4453 -10960 4853 -10922
rect 4453 -10994 4469 -10960
rect 4837 -10994 4853 -10960
rect 4453 -11010 4853 -10994
rect 5373 -10960 5773 -10922
rect 5373 -10994 5389 -10960
rect 5757 -10994 5773 -10960
rect 5373 -11010 5773 -10994
rect 6376 -10130 6576 -10114
rect 6376 -10164 6392 -10130
rect 6560 -10164 6576 -10130
rect 6376 -10211 6576 -10164
rect 6376 -10358 6576 -10311
rect 6376 -10392 6392 -10358
rect 6560 -10392 6576 -10358
rect 6376 -10408 6576 -10392
rect 6376 -10698 6576 -10682
rect 6376 -10732 6392 -10698
rect 6560 -10732 6576 -10698
rect 6376 -10770 6576 -10732
rect 6376 -10908 6576 -10870
rect 6376 -10942 6392 -10908
rect 6560 -10942 6576 -10908
rect 6376 -10958 6576 -10942
<< polycont >>
rect -1127 2592 -1093 2626
rect -1029 2592 -995 2626
rect -931 2592 -897 2626
rect -833 2592 -799 2626
rect -735 2592 -701 2626
rect -637 2592 -603 2626
rect -539 2592 -505 2626
rect -441 2592 -407 2626
rect -343 2592 -309 2626
rect -245 2592 -211 2626
rect -147 2592 -113 2626
rect -49 2592 -15 2626
rect 49 2592 83 2626
rect 147 2592 181 2626
rect 245 2592 279 2626
rect -1127 2064 -1093 2098
rect -1029 2064 -995 2098
rect -931 2064 -897 2098
rect -833 2064 -799 2098
rect -735 2064 -701 2098
rect -637 2064 -603 2098
rect -539 2064 -505 2098
rect -441 2064 -407 2098
rect -343 2064 -309 2098
rect -245 2064 -211 2098
rect -147 2064 -113 2098
rect -49 2064 -15 2098
rect 49 2064 83 2098
rect 147 2064 181 2098
rect 245 2064 279 2098
rect -1127 1956 -1093 1990
rect -1029 1956 -995 1990
rect -931 1956 -897 1990
rect -833 1956 -799 1990
rect -735 1956 -701 1990
rect -637 1956 -603 1990
rect -539 1956 -505 1990
rect -441 1956 -407 1990
rect -343 1956 -309 1990
rect -245 1956 -211 1990
rect -147 1956 -113 1990
rect -49 1956 -15 1990
rect 49 1956 83 1990
rect 147 1956 181 1990
rect 245 1956 279 1990
rect -1127 1428 -1093 1462
rect -1029 1428 -995 1462
rect -931 1428 -897 1462
rect -833 1428 -799 1462
rect -735 1428 -701 1462
rect -637 1428 -603 1462
rect -539 1428 -505 1462
rect -441 1428 -407 1462
rect -343 1428 -309 1462
rect -245 1428 -211 1462
rect -147 1428 -113 1462
rect -49 1428 -15 1462
rect 49 1428 83 1462
rect 147 1428 181 1462
rect 245 1428 279 1462
rect 671 2592 705 2626
rect 769 2592 803 2626
rect 867 2592 901 2626
rect 965 2592 999 2626
rect 1063 2592 1097 2626
rect 1161 2592 1195 2626
rect 1259 2592 1293 2626
rect 1357 2592 1391 2626
rect 1455 2592 1489 2626
rect 1553 2592 1587 2626
rect 1651 2592 1685 2626
rect 1749 2592 1783 2626
rect 1847 2592 1881 2626
rect 1945 2592 1979 2626
rect 2043 2592 2077 2626
rect 671 2064 705 2098
rect 769 2064 803 2098
rect 867 2064 901 2098
rect 965 2064 999 2098
rect 1063 2064 1097 2098
rect 1161 2064 1195 2098
rect 1259 2064 1293 2098
rect 1357 2064 1391 2098
rect 1455 2064 1489 2098
rect 1553 2064 1587 2098
rect 1651 2064 1685 2098
rect 1749 2064 1783 2098
rect 1847 2064 1881 2098
rect 1945 2064 1979 2098
rect 2043 2064 2077 2098
rect 671 1956 705 1990
rect 769 1956 803 1990
rect 867 1956 901 1990
rect 965 1956 999 1990
rect 1063 1956 1097 1990
rect 1161 1956 1195 1990
rect 1259 1956 1293 1990
rect 1357 1956 1391 1990
rect 1455 1956 1489 1990
rect 1553 1956 1587 1990
rect 1651 1956 1685 1990
rect 1749 1956 1783 1990
rect 1847 1956 1881 1990
rect 1945 1956 1979 1990
rect 2043 1956 2077 1990
rect 671 1428 705 1462
rect 769 1428 803 1462
rect 867 1428 901 1462
rect 965 1428 999 1462
rect 1063 1428 1097 1462
rect 1161 1428 1195 1462
rect 1259 1428 1293 1462
rect 1357 1428 1391 1462
rect 1455 1428 1489 1462
rect 1553 1428 1587 1462
rect 1651 1428 1685 1462
rect 1749 1428 1783 1462
rect 1847 1428 1881 1462
rect 1945 1428 1979 1462
rect 2043 1428 2077 1462
rect 2486 1940 2554 1974
rect 2644 1940 2712 1974
rect 2802 1940 2870 1974
rect 2960 1940 3028 1974
rect 3118 1940 3186 1974
rect 3276 1940 3344 1974
rect 3434 1940 3502 1974
rect 3592 1940 3660 1974
rect 3750 1940 3818 1974
rect 3908 1940 3976 1974
rect 2486 1412 2554 1446
rect 2644 1412 2712 1446
rect 2802 1412 2870 1446
rect 2960 1412 3028 1446
rect 3118 1412 3186 1446
rect 3276 1412 3344 1446
rect 3434 1412 3502 1446
rect 3592 1412 3660 1446
rect 3750 1412 3818 1446
rect 3908 1412 3976 1446
rect -1127 1116 -1093 1150
rect -1030 1116 -996 1150
rect -931 1116 -897 1150
rect -834 1116 -800 1150
rect -735 1116 -701 1150
rect -638 1116 -604 1150
rect -539 1116 -505 1150
rect -442 1116 -408 1150
rect -343 1116 -309 1150
rect -246 1116 -212 1150
rect -147 1116 -113 1150
rect -50 1116 -16 1150
rect 49 1116 83 1150
rect 146 1116 180 1150
rect 245 1116 279 1150
rect 342 1116 376 1150
rect 441 1116 475 1150
rect 538 1116 572 1150
rect 637 1116 671 1150
rect 734 1116 768 1150
rect 833 1116 867 1150
rect 930 1116 964 1150
rect 1029 1116 1063 1150
rect 1126 1116 1160 1150
rect 1225 1116 1259 1150
rect -1128 606 -1094 640
rect -1029 606 -995 640
rect -932 606 -898 640
rect -833 606 -799 640
rect -736 606 -702 640
rect -637 606 -603 640
rect -540 606 -506 640
rect -441 606 -407 640
rect -344 606 -310 640
rect -245 606 -211 640
rect -148 606 -114 640
rect -49 606 -15 640
rect 48 606 82 640
rect 147 606 181 640
rect 244 606 278 640
rect 343 606 377 640
rect 440 606 474 640
rect 539 606 573 640
rect 636 606 670 640
rect 735 606 769 640
rect 832 606 866 640
rect 931 606 965 640
rect 1028 606 1062 640
rect 1127 606 1161 640
rect 1224 606 1258 640
rect -1127 498 -1093 532
rect -1029 498 -995 532
rect -931 498 -897 532
rect -833 498 -799 532
rect -735 498 -701 532
rect -637 498 -603 532
rect -539 498 -505 532
rect -441 498 -407 532
rect -343 498 -309 532
rect -245 498 -211 532
rect -147 498 -113 532
rect -49 498 -15 532
rect 49 498 83 532
rect 147 498 181 532
rect 245 498 279 532
rect 343 498 377 532
rect 441 498 475 532
rect 539 498 573 532
rect 637 498 671 532
rect 735 498 769 532
rect 833 498 867 532
rect 931 498 965 532
rect 1029 498 1063 532
rect 1127 498 1161 532
rect 1225 498 1259 532
rect -1127 -12 -1093 22
rect -1029 -12 -995 22
rect -931 -12 -897 22
rect -833 -12 -799 22
rect -735 -12 -701 22
rect -637 -12 -603 22
rect -539 -12 -505 22
rect -441 -12 -407 22
rect -343 -12 -309 22
rect -245 -12 -211 22
rect -147 -12 -113 22
rect -49 -12 -15 22
rect 49 -12 83 22
rect 147 -12 181 22
rect 245 -12 279 22
rect 343 -12 377 22
rect 441 -12 475 22
rect 539 -12 573 22
rect 637 -12 671 22
rect 735 -12 769 22
rect 833 -12 867 22
rect 931 -12 965 22
rect 1029 -12 1063 22
rect 1127 -12 1161 22
rect 1225 -12 1259 22
rect -1127 -328 -1093 -294
rect -1030 -328 -996 -294
rect -931 -328 -897 -294
rect -834 -328 -800 -294
rect -735 -328 -701 -294
rect -638 -328 -604 -294
rect -539 -328 -505 -294
rect -442 -328 -408 -294
rect -343 -328 -309 -294
rect -246 -328 -212 -294
rect -147 -328 -113 -294
rect -50 -328 -16 -294
rect 49 -328 83 -294
rect 146 -328 180 -294
rect 245 -328 279 -294
rect 342 -328 376 -294
rect 441 -328 475 -294
rect 538 -328 572 -294
rect 637 -328 671 -294
rect 734 -328 768 -294
rect 833 -328 867 -294
rect 930 -328 964 -294
rect 1029 -328 1063 -294
rect 1126 -328 1160 -294
rect 1225 -328 1259 -294
rect -1128 -838 -1094 -804
rect -1029 -838 -995 -804
rect -932 -838 -898 -804
rect -833 -838 -799 -804
rect -736 -838 -702 -804
rect -637 -838 -603 -804
rect -540 -838 -506 -804
rect -441 -838 -407 -804
rect -344 -838 -310 -804
rect -245 -838 -211 -804
rect -148 -838 -114 -804
rect -49 -838 -15 -804
rect 48 -838 82 -804
rect 147 -838 181 -804
rect 244 -838 278 -804
rect 343 -838 377 -804
rect 440 -838 474 -804
rect 539 -838 573 -804
rect 636 -838 670 -804
rect 735 -838 769 -804
rect 832 -838 866 -804
rect 931 -838 965 -804
rect 1028 -838 1062 -804
rect 1127 -838 1161 -804
rect 1224 -838 1258 -804
rect -1127 -946 -1093 -912
rect -1029 -946 -995 -912
rect -931 -946 -897 -912
rect -833 -946 -799 -912
rect -735 -946 -701 -912
rect -637 -946 -603 -912
rect -539 -946 -505 -912
rect -441 -946 -407 -912
rect -343 -946 -309 -912
rect -245 -946 -211 -912
rect -147 -946 -113 -912
rect -49 -946 -15 -912
rect 49 -946 83 -912
rect 147 -946 181 -912
rect 245 -946 279 -912
rect 343 -946 377 -912
rect 441 -946 475 -912
rect 539 -946 573 -912
rect 637 -946 671 -912
rect 735 -946 769 -912
rect 833 -946 867 -912
rect 931 -946 965 -912
rect 1029 -946 1063 -912
rect 1127 -946 1161 -912
rect 1225 -946 1259 -912
rect -1127 -1456 -1093 -1422
rect -1029 -1456 -995 -1422
rect -931 -1456 -897 -1422
rect -833 -1456 -799 -1422
rect -735 -1456 -701 -1422
rect -637 -1456 -603 -1422
rect -539 -1456 -505 -1422
rect -441 -1456 -407 -1422
rect -343 -1456 -309 -1422
rect -245 -1456 -211 -1422
rect -147 -1456 -113 -1422
rect -49 -1456 -15 -1422
rect 49 -1456 83 -1422
rect 147 -1456 181 -1422
rect 245 -1456 279 -1422
rect 343 -1456 377 -1422
rect 441 -1456 475 -1422
rect 539 -1456 573 -1422
rect 637 -1456 671 -1422
rect 735 -1456 769 -1422
rect 833 -1456 867 -1422
rect 931 -1456 965 -1422
rect 1029 -1456 1063 -1422
rect 1127 -1456 1161 -1422
rect 1225 -1456 1259 -1422
rect 2533 796 2567 830
rect 2631 796 2665 830
rect 2729 796 2763 830
rect 2827 796 2861 830
rect 2925 796 2959 830
rect 3023 796 3057 830
rect 3121 796 3155 830
rect 3219 796 3253 830
rect 3317 796 3351 830
rect 3415 796 3449 830
rect 3513 796 3547 830
rect 3611 796 3645 830
rect 3709 796 3743 830
rect 3807 796 3841 830
rect 3905 796 3939 830
rect 2533 286 2567 320
rect 2631 286 2665 320
rect 2729 286 2763 320
rect 2827 286 2861 320
rect 2925 286 2959 320
rect 3023 286 3057 320
rect 3121 286 3155 320
rect 3219 286 3253 320
rect 3317 286 3351 320
rect 3415 286 3449 320
rect 3513 286 3547 320
rect 3611 286 3645 320
rect 3709 286 3743 320
rect 3807 286 3841 320
rect 3905 286 3939 320
rect 2533 178 2567 212
rect 2631 178 2665 212
rect 2729 178 2763 212
rect 2827 178 2861 212
rect 2925 178 2959 212
rect 3023 178 3057 212
rect 3121 178 3155 212
rect 3219 178 3253 212
rect 3317 178 3351 212
rect 3415 178 3449 212
rect 3513 178 3547 212
rect 3611 178 3645 212
rect 3709 178 3743 212
rect 3807 178 3841 212
rect 3905 178 3939 212
rect 2533 -332 2567 -298
rect 2631 -332 2665 -298
rect 2729 -332 2763 -298
rect 2827 -332 2861 -298
rect 2925 -332 2959 -298
rect 3023 -332 3057 -298
rect 3121 -332 3155 -298
rect 3219 -332 3253 -298
rect 3317 -332 3351 -298
rect 3415 -332 3449 -298
rect 3513 -332 3547 -298
rect 3611 -332 3645 -298
rect 3709 -332 3743 -298
rect 3807 -332 3841 -298
rect 3905 -332 3939 -298
rect 1662 -982 1696 -948
rect 1758 -982 1792 -948
rect 1854 -982 1888 -948
rect 1950 -982 1984 -948
rect 2046 -982 2080 -948
rect 2142 -982 2176 -948
rect 2238 -982 2272 -948
rect 2334 -982 2368 -948
rect 2430 -982 2464 -948
rect 2526 -982 2560 -948
rect 2622 -982 2656 -948
rect 2718 -982 2752 -948
rect 1662 -1492 1696 -1458
rect 1758 -1492 1792 -1458
rect 1854 -1492 1888 -1458
rect 1950 -1492 1984 -1458
rect 2046 -1492 2080 -1458
rect 2142 -1492 2176 -1458
rect 2238 -1492 2272 -1458
rect 2334 -1492 2368 -1458
rect 2430 -1492 2464 -1458
rect 2526 -1492 2560 -1458
rect 2622 -1492 2656 -1458
rect 2718 -1492 2752 -1458
rect -1148 -1748 -1114 -1714
rect -956 -1748 -922 -1714
rect -764 -1748 -730 -1714
rect -572 -1748 -538 -1714
rect -380 -1748 -346 -1714
rect -188 -1748 -154 -1714
rect 4 -1748 38 -1714
rect 196 -1748 230 -1714
rect 388 -1748 422 -1714
rect 580 -1748 614 -1714
rect 772 -1748 806 -1714
rect 964 -1748 998 -1714
rect 1156 -1748 1190 -1714
rect -1052 -2258 -1018 -2224
rect -860 -2258 -826 -2224
rect -668 -2258 -634 -2224
rect -476 -2258 -442 -2224
rect -284 -2258 -250 -2224
rect -92 -2258 -58 -2224
rect 100 -2258 134 -2224
rect 292 -2258 326 -2224
rect 484 -2258 518 -2224
rect 676 -2258 710 -2224
rect 868 -2258 902 -2224
rect 1060 -2258 1094 -2224
rect -1052 -2366 -1018 -2332
rect -860 -2366 -826 -2332
rect -668 -2366 -634 -2332
rect -476 -2366 -442 -2332
rect -284 -2366 -250 -2332
rect -92 -2366 -58 -2332
rect 100 -2366 134 -2332
rect 292 -2366 326 -2332
rect 484 -2366 518 -2332
rect 676 -2366 710 -2332
rect 868 -2366 902 -2332
rect 1060 -2366 1094 -2332
rect -1148 -2876 -1114 -2842
rect -956 -2876 -922 -2842
rect -764 -2876 -730 -2842
rect -572 -2876 -538 -2842
rect -380 -2876 -346 -2842
rect -188 -2876 -154 -2842
rect 4 -2876 38 -2842
rect 196 -2876 230 -2842
rect 388 -2876 422 -2842
rect 580 -2876 614 -2842
rect 772 -2876 806 -2842
rect 964 -2876 998 -2842
rect 1156 -2876 1190 -2842
rect -1148 -2984 -1114 -2950
rect -956 -2984 -922 -2950
rect -764 -2984 -730 -2950
rect -572 -2984 -538 -2950
rect -380 -2984 -346 -2950
rect -188 -2984 -154 -2950
rect 4 -2984 38 -2950
rect 196 -2984 230 -2950
rect 388 -2984 422 -2950
rect 580 -2984 614 -2950
rect 772 -2984 806 -2950
rect 964 -2984 998 -2950
rect 1156 -2984 1190 -2950
rect -1052 -3494 -1018 -3460
rect -860 -3494 -826 -3460
rect -668 -3494 -634 -3460
rect -476 -3494 -442 -3460
rect -284 -3494 -250 -3460
rect -92 -3494 -58 -3460
rect 100 -3494 134 -3460
rect 292 -3494 326 -3460
rect 484 -3494 518 -3460
rect 676 -3494 710 -3460
rect 868 -3494 902 -3460
rect 1060 -3494 1094 -3460
rect -1052 -3602 -1018 -3568
rect -860 -3602 -826 -3568
rect -668 -3602 -634 -3568
rect -476 -3602 -442 -3568
rect -284 -3602 -250 -3568
rect -92 -3602 -58 -3568
rect 100 -3602 134 -3568
rect 292 -3602 326 -3568
rect 484 -3602 518 -3568
rect 676 -3602 710 -3568
rect 868 -3602 902 -3568
rect 1060 -3602 1094 -3568
rect -1148 -4112 -1114 -4078
rect -956 -4112 -922 -4078
rect -764 -4112 -730 -4078
rect -572 -4112 -538 -4078
rect -380 -4112 -346 -4078
rect -188 -4112 -154 -4078
rect 4 -4112 38 -4078
rect 196 -4112 230 -4078
rect 388 -4112 422 -4078
rect 580 -4112 614 -4078
rect 772 -4112 806 -4078
rect 964 -4112 998 -4078
rect 1156 -4112 1190 -4078
rect 1676 -1802 1844 -1768
rect 1934 -1802 2102 -1768
rect 2192 -1802 2360 -1768
rect 2450 -1802 2618 -1768
rect 2708 -1802 2876 -1768
rect 2966 -1802 3134 -1768
rect 1676 -2312 1844 -2278
rect 1934 -2312 2102 -2278
rect 2192 -2312 2360 -2278
rect 2450 -2312 2618 -2278
rect 2708 -2312 2876 -2278
rect 2966 -2312 3134 -2278
rect -1127 -4478 -1093 -4444
rect -1029 -4478 -995 -4444
rect -931 -4478 -897 -4444
rect -833 -4478 -799 -4444
rect -735 -4478 -701 -4444
rect -637 -4478 -603 -4444
rect -539 -4478 -505 -4444
rect -441 -4478 -407 -4444
rect -343 -4478 -309 -4444
rect -245 -4478 -211 -4444
rect -147 -4478 -113 -4444
rect -49 -4478 -15 -4444
rect 49 -4478 83 -4444
rect 147 -4478 181 -4444
rect 245 -4478 279 -4444
rect -1127 -5006 -1093 -4972
rect -1029 -5006 -995 -4972
rect -931 -5006 -897 -4972
rect -833 -5006 -799 -4972
rect -735 -5006 -701 -4972
rect -637 -5006 -603 -4972
rect -539 -5006 -505 -4972
rect -441 -5006 -407 -4972
rect -343 -5006 -309 -4972
rect -245 -5006 -211 -4972
rect -147 -5006 -113 -4972
rect -49 -5006 -15 -4972
rect 49 -5006 83 -4972
rect 147 -5006 181 -4972
rect 245 -5006 279 -4972
rect -1127 -5114 -1093 -5080
rect -1029 -5114 -995 -5080
rect -931 -5114 -897 -5080
rect -833 -5114 -799 -5080
rect -735 -5114 -701 -5080
rect -637 -5114 -603 -5080
rect -539 -5114 -505 -5080
rect -441 -5114 -407 -5080
rect -343 -5114 -309 -5080
rect -245 -5114 -211 -5080
rect -147 -5114 -113 -5080
rect -49 -5114 -15 -5080
rect 49 -5114 83 -5080
rect 147 -5114 181 -5080
rect 245 -5114 279 -5080
rect -1127 -5642 -1093 -5608
rect -1029 -5642 -995 -5608
rect -931 -5642 -897 -5608
rect -833 -5642 -799 -5608
rect -735 -5642 -701 -5608
rect -637 -5642 -603 -5608
rect -539 -5642 -505 -5608
rect -441 -5642 -407 -5608
rect -343 -5642 -309 -5608
rect -245 -5642 -211 -5608
rect -147 -5642 -113 -5608
rect -49 -5642 -15 -5608
rect 49 -5642 83 -5608
rect 147 -5642 181 -5608
rect 245 -5642 279 -5608
rect 671 -4478 705 -4444
rect 769 -4478 803 -4444
rect 867 -4478 901 -4444
rect 965 -4478 999 -4444
rect 1063 -4478 1097 -4444
rect 1161 -4478 1195 -4444
rect 1259 -4478 1293 -4444
rect 1357 -4478 1391 -4444
rect 1455 -4478 1489 -4444
rect 1553 -4478 1587 -4444
rect 1651 -4478 1685 -4444
rect 1749 -4478 1783 -4444
rect 1847 -4478 1881 -4444
rect 1945 -4478 1979 -4444
rect 2043 -4478 2077 -4444
rect 671 -5006 705 -4972
rect 769 -5006 803 -4972
rect 867 -5006 901 -4972
rect 965 -5006 999 -4972
rect 1063 -5006 1097 -4972
rect 1161 -5006 1195 -4972
rect 1259 -5006 1293 -4972
rect 1357 -5006 1391 -4972
rect 1455 -5006 1489 -4972
rect 1553 -5006 1587 -4972
rect 1651 -5006 1685 -4972
rect 1749 -5006 1783 -4972
rect 1847 -5006 1881 -4972
rect 1945 -5006 1979 -4972
rect 2043 -5006 2077 -4972
rect 671 -5114 705 -5080
rect 769 -5114 803 -5080
rect 867 -5114 901 -5080
rect 965 -5114 999 -5080
rect 1063 -5114 1097 -5080
rect 1161 -5114 1195 -5080
rect 1259 -5114 1293 -5080
rect 1357 -5114 1391 -5080
rect 1455 -5114 1489 -5080
rect 1553 -5114 1587 -5080
rect 1651 -5114 1685 -5080
rect 1749 -5114 1783 -5080
rect 1847 -5114 1881 -5080
rect 1945 -5114 1979 -5080
rect 2043 -5114 2077 -5080
rect 671 -5642 705 -5608
rect 769 -5642 803 -5608
rect 867 -5642 901 -5608
rect 965 -5642 999 -5608
rect 1063 -5642 1097 -5608
rect 1161 -5642 1195 -5608
rect 1259 -5642 1293 -5608
rect 1357 -5642 1391 -5608
rect 1455 -5642 1489 -5608
rect 1553 -5642 1587 -5608
rect 1651 -5642 1685 -5608
rect 1749 -5642 1783 -5608
rect 1847 -5642 1881 -5608
rect 1945 -5642 1979 -5608
rect 2043 -5642 2077 -5608
rect 2486 -5130 2554 -5096
rect 2644 -5130 2712 -5096
rect 2802 -5130 2870 -5096
rect 2960 -5130 3028 -5096
rect 3118 -5130 3186 -5096
rect 3276 -5130 3344 -5096
rect 3434 -5130 3502 -5096
rect 3592 -5130 3660 -5096
rect 3750 -5130 3818 -5096
rect 3908 -5130 3976 -5096
rect 2486 -5658 2554 -5624
rect 2644 -5658 2712 -5624
rect 2802 -5658 2870 -5624
rect 2960 -5658 3028 -5624
rect 3118 -5658 3186 -5624
rect 3276 -5658 3344 -5624
rect 3434 -5658 3502 -5624
rect 3592 -5658 3660 -5624
rect 3750 -5658 3818 -5624
rect 3908 -5658 3976 -5624
rect -1127 -5954 -1093 -5920
rect -1030 -5954 -996 -5920
rect -931 -5954 -897 -5920
rect -834 -5954 -800 -5920
rect -735 -5954 -701 -5920
rect -638 -5954 -604 -5920
rect -539 -5954 -505 -5920
rect -442 -5954 -408 -5920
rect -343 -5954 -309 -5920
rect -246 -5954 -212 -5920
rect -147 -5954 -113 -5920
rect -50 -5954 -16 -5920
rect 49 -5954 83 -5920
rect 146 -5954 180 -5920
rect 245 -5954 279 -5920
rect 342 -5954 376 -5920
rect 441 -5954 475 -5920
rect 538 -5954 572 -5920
rect 637 -5954 671 -5920
rect 734 -5954 768 -5920
rect 833 -5954 867 -5920
rect 930 -5954 964 -5920
rect 1029 -5954 1063 -5920
rect 1126 -5954 1160 -5920
rect 1225 -5954 1259 -5920
rect -1128 -6464 -1094 -6430
rect -1029 -6464 -995 -6430
rect -932 -6464 -898 -6430
rect -833 -6464 -799 -6430
rect -736 -6464 -702 -6430
rect -637 -6464 -603 -6430
rect -540 -6464 -506 -6430
rect -441 -6464 -407 -6430
rect -344 -6464 -310 -6430
rect -245 -6464 -211 -6430
rect -148 -6464 -114 -6430
rect -49 -6464 -15 -6430
rect 48 -6464 82 -6430
rect 147 -6464 181 -6430
rect 244 -6464 278 -6430
rect 343 -6464 377 -6430
rect 440 -6464 474 -6430
rect 539 -6464 573 -6430
rect 636 -6464 670 -6430
rect 735 -6464 769 -6430
rect 832 -6464 866 -6430
rect 931 -6464 965 -6430
rect 1028 -6464 1062 -6430
rect 1127 -6464 1161 -6430
rect 1224 -6464 1258 -6430
rect -1127 -6572 -1093 -6538
rect -1029 -6572 -995 -6538
rect -931 -6572 -897 -6538
rect -833 -6572 -799 -6538
rect -735 -6572 -701 -6538
rect -637 -6572 -603 -6538
rect -539 -6572 -505 -6538
rect -441 -6572 -407 -6538
rect -343 -6572 -309 -6538
rect -245 -6572 -211 -6538
rect -147 -6572 -113 -6538
rect -49 -6572 -15 -6538
rect 49 -6572 83 -6538
rect 147 -6572 181 -6538
rect 245 -6572 279 -6538
rect 343 -6572 377 -6538
rect 441 -6572 475 -6538
rect 539 -6572 573 -6538
rect 637 -6572 671 -6538
rect 735 -6572 769 -6538
rect 833 -6572 867 -6538
rect 931 -6572 965 -6538
rect 1029 -6572 1063 -6538
rect 1127 -6572 1161 -6538
rect 1225 -6572 1259 -6538
rect -1127 -7082 -1093 -7048
rect -1029 -7082 -995 -7048
rect -931 -7082 -897 -7048
rect -833 -7082 -799 -7048
rect -735 -7082 -701 -7048
rect -637 -7082 -603 -7048
rect -539 -7082 -505 -7048
rect -441 -7082 -407 -7048
rect -343 -7082 -309 -7048
rect -245 -7082 -211 -7048
rect -147 -7082 -113 -7048
rect -49 -7082 -15 -7048
rect 49 -7082 83 -7048
rect 147 -7082 181 -7048
rect 245 -7082 279 -7048
rect 343 -7082 377 -7048
rect 441 -7082 475 -7048
rect 539 -7082 573 -7048
rect 637 -7082 671 -7048
rect 735 -7082 769 -7048
rect 833 -7082 867 -7048
rect 931 -7082 965 -7048
rect 1029 -7082 1063 -7048
rect 1127 -7082 1161 -7048
rect 1225 -7082 1259 -7048
rect -1127 -7398 -1093 -7364
rect -1030 -7398 -996 -7364
rect -931 -7398 -897 -7364
rect -834 -7398 -800 -7364
rect -735 -7398 -701 -7364
rect -638 -7398 -604 -7364
rect -539 -7398 -505 -7364
rect -442 -7398 -408 -7364
rect -343 -7398 -309 -7364
rect -246 -7398 -212 -7364
rect -147 -7398 -113 -7364
rect -50 -7398 -16 -7364
rect 49 -7398 83 -7364
rect 146 -7398 180 -7364
rect 245 -7398 279 -7364
rect 342 -7398 376 -7364
rect 441 -7398 475 -7364
rect 538 -7398 572 -7364
rect 637 -7398 671 -7364
rect 734 -7398 768 -7364
rect 833 -7398 867 -7364
rect 930 -7398 964 -7364
rect 1029 -7398 1063 -7364
rect 1126 -7398 1160 -7364
rect 1225 -7398 1259 -7364
rect -1128 -7908 -1094 -7874
rect -1029 -7908 -995 -7874
rect -932 -7908 -898 -7874
rect -833 -7908 -799 -7874
rect -736 -7908 -702 -7874
rect -637 -7908 -603 -7874
rect -540 -7908 -506 -7874
rect -441 -7908 -407 -7874
rect -344 -7908 -310 -7874
rect -245 -7908 -211 -7874
rect -148 -7908 -114 -7874
rect -49 -7908 -15 -7874
rect 48 -7908 82 -7874
rect 147 -7908 181 -7874
rect 244 -7908 278 -7874
rect 343 -7908 377 -7874
rect 440 -7908 474 -7874
rect 539 -7908 573 -7874
rect 636 -7908 670 -7874
rect 735 -7908 769 -7874
rect 832 -7908 866 -7874
rect 931 -7908 965 -7874
rect 1028 -7908 1062 -7874
rect 1127 -7908 1161 -7874
rect 1224 -7908 1258 -7874
rect -1127 -8016 -1093 -7982
rect -1029 -8016 -995 -7982
rect -931 -8016 -897 -7982
rect -833 -8016 -799 -7982
rect -735 -8016 -701 -7982
rect -637 -8016 -603 -7982
rect -539 -8016 -505 -7982
rect -441 -8016 -407 -7982
rect -343 -8016 -309 -7982
rect -245 -8016 -211 -7982
rect -147 -8016 -113 -7982
rect -49 -8016 -15 -7982
rect 49 -8016 83 -7982
rect 147 -8016 181 -7982
rect 245 -8016 279 -7982
rect 343 -8016 377 -7982
rect 441 -8016 475 -7982
rect 539 -8016 573 -7982
rect 637 -8016 671 -7982
rect 735 -8016 769 -7982
rect 833 -8016 867 -7982
rect 931 -8016 965 -7982
rect 1029 -8016 1063 -7982
rect 1127 -8016 1161 -7982
rect 1225 -8016 1259 -7982
rect -1127 -8526 -1093 -8492
rect -1029 -8526 -995 -8492
rect -931 -8526 -897 -8492
rect -833 -8526 -799 -8492
rect -735 -8526 -701 -8492
rect -637 -8526 -603 -8492
rect -539 -8526 -505 -8492
rect -441 -8526 -407 -8492
rect -343 -8526 -309 -8492
rect -245 -8526 -211 -8492
rect -147 -8526 -113 -8492
rect -49 -8526 -15 -8492
rect 49 -8526 83 -8492
rect 147 -8526 181 -8492
rect 245 -8526 279 -8492
rect 343 -8526 377 -8492
rect 441 -8526 475 -8492
rect 539 -8526 573 -8492
rect 637 -8526 671 -8492
rect 735 -8526 769 -8492
rect 833 -8526 867 -8492
rect 931 -8526 965 -8492
rect 1029 -8526 1063 -8492
rect 1127 -8526 1161 -8492
rect 1225 -8526 1259 -8492
rect 2533 -6274 2567 -6240
rect 2631 -6274 2665 -6240
rect 2729 -6274 2763 -6240
rect 2827 -6274 2861 -6240
rect 2925 -6274 2959 -6240
rect 3023 -6274 3057 -6240
rect 3121 -6274 3155 -6240
rect 3219 -6274 3253 -6240
rect 3317 -6274 3351 -6240
rect 3415 -6274 3449 -6240
rect 3513 -6274 3547 -6240
rect 3611 -6274 3645 -6240
rect 3709 -6274 3743 -6240
rect 3807 -6274 3841 -6240
rect 3905 -6274 3939 -6240
rect 2533 -6784 2567 -6750
rect 2631 -6784 2665 -6750
rect 2729 -6784 2763 -6750
rect 2827 -6784 2861 -6750
rect 2925 -6784 2959 -6750
rect 3023 -6784 3057 -6750
rect 3121 -6784 3155 -6750
rect 3219 -6784 3253 -6750
rect 3317 -6784 3351 -6750
rect 3415 -6784 3449 -6750
rect 3513 -6784 3547 -6750
rect 3611 -6784 3645 -6750
rect 3709 -6784 3743 -6750
rect 3807 -6784 3841 -6750
rect 3905 -6784 3939 -6750
rect 2533 -6892 2567 -6858
rect 2631 -6892 2665 -6858
rect 2729 -6892 2763 -6858
rect 2827 -6892 2861 -6858
rect 2925 -6892 2959 -6858
rect 3023 -6892 3057 -6858
rect 3121 -6892 3155 -6858
rect 3219 -6892 3253 -6858
rect 3317 -6892 3351 -6858
rect 3415 -6892 3449 -6858
rect 3513 -6892 3547 -6858
rect 3611 -6892 3645 -6858
rect 3709 -6892 3743 -6858
rect 3807 -6892 3841 -6858
rect 3905 -6892 3939 -6858
rect 2533 -7402 2567 -7368
rect 2631 -7402 2665 -7368
rect 2729 -7402 2763 -7368
rect 2827 -7402 2861 -7368
rect 2925 -7402 2959 -7368
rect 3023 -7402 3057 -7368
rect 3121 -7402 3155 -7368
rect 3219 -7402 3253 -7368
rect 3317 -7402 3351 -7368
rect 3415 -7402 3449 -7368
rect 3513 -7402 3547 -7368
rect 3611 -7402 3645 -7368
rect 3709 -7402 3743 -7368
rect 3807 -7402 3841 -7368
rect 3905 -7402 3939 -7368
rect 1662 -8052 1696 -8018
rect 1758 -8052 1792 -8018
rect 1854 -8052 1888 -8018
rect 1950 -8052 1984 -8018
rect 2046 -8052 2080 -8018
rect 2142 -8052 2176 -8018
rect 2238 -8052 2272 -8018
rect 2334 -8052 2368 -8018
rect 2430 -8052 2464 -8018
rect 2526 -8052 2560 -8018
rect 2622 -8052 2656 -8018
rect 2718 -8052 2752 -8018
rect 1662 -8562 1696 -8528
rect 1758 -8562 1792 -8528
rect 1854 -8562 1888 -8528
rect 1950 -8562 1984 -8528
rect 2046 -8562 2080 -8528
rect 2142 -8562 2176 -8528
rect 2238 -8562 2272 -8528
rect 2334 -8562 2368 -8528
rect 2430 -8562 2464 -8528
rect 2526 -8562 2560 -8528
rect 2622 -8562 2656 -8528
rect 2718 -8562 2752 -8528
rect 3558 -8052 3592 -8018
rect 3654 -8052 3688 -8018
rect 3750 -8052 3784 -8018
rect 3846 -8052 3880 -8018
rect 3942 -8052 3976 -8018
rect 4038 -8052 4072 -8018
rect 4134 -8052 4168 -8018
rect 4230 -8052 4264 -8018
rect 4326 -8052 4360 -8018
rect 4422 -8052 4456 -8018
rect 4518 -8052 4552 -8018
rect 4614 -8052 4648 -8018
rect 3558 -8562 3592 -8528
rect 3654 -8562 3688 -8528
rect 3750 -8562 3784 -8528
rect 3846 -8562 3880 -8528
rect 3942 -8562 3976 -8528
rect 4038 -8562 4072 -8528
rect 4134 -8562 4168 -8528
rect 4230 -8562 4264 -8528
rect 4326 -8562 4360 -8528
rect 4422 -8562 4456 -8528
rect 4518 -8562 4552 -8528
rect 4614 -8562 4648 -8528
rect -1148 -8818 -1114 -8784
rect -956 -8818 -922 -8784
rect -764 -8818 -730 -8784
rect -572 -8818 -538 -8784
rect -380 -8818 -346 -8784
rect -188 -8818 -154 -8784
rect 4 -8818 38 -8784
rect 196 -8818 230 -8784
rect 388 -8818 422 -8784
rect 580 -8818 614 -8784
rect 772 -8818 806 -8784
rect 964 -8818 998 -8784
rect 1156 -8818 1190 -8784
rect -1052 -9328 -1018 -9294
rect -860 -9328 -826 -9294
rect -668 -9328 -634 -9294
rect -476 -9328 -442 -9294
rect -284 -9328 -250 -9294
rect -92 -9328 -58 -9294
rect 100 -9328 134 -9294
rect 292 -9328 326 -9294
rect 484 -9328 518 -9294
rect 676 -9328 710 -9294
rect 868 -9328 902 -9294
rect 1060 -9328 1094 -9294
rect -1052 -9436 -1018 -9402
rect -860 -9436 -826 -9402
rect -668 -9436 -634 -9402
rect -476 -9436 -442 -9402
rect -284 -9436 -250 -9402
rect -92 -9436 -58 -9402
rect 100 -9436 134 -9402
rect 292 -9436 326 -9402
rect 484 -9436 518 -9402
rect 676 -9436 710 -9402
rect 868 -9436 902 -9402
rect 1060 -9436 1094 -9402
rect -1148 -9946 -1114 -9912
rect -956 -9946 -922 -9912
rect -764 -9946 -730 -9912
rect -572 -9946 -538 -9912
rect -380 -9946 -346 -9912
rect -188 -9946 -154 -9912
rect 4 -9946 38 -9912
rect 196 -9946 230 -9912
rect 388 -9946 422 -9912
rect 580 -9946 614 -9912
rect 772 -9946 806 -9912
rect 964 -9946 998 -9912
rect 1156 -9946 1190 -9912
rect -1148 -10054 -1114 -10020
rect -956 -10054 -922 -10020
rect -764 -10054 -730 -10020
rect -572 -10054 -538 -10020
rect -380 -10054 -346 -10020
rect -188 -10054 -154 -10020
rect 4 -10054 38 -10020
rect 196 -10054 230 -10020
rect 388 -10054 422 -10020
rect 580 -10054 614 -10020
rect 772 -10054 806 -10020
rect 964 -10054 998 -10020
rect 1156 -10054 1190 -10020
rect -1052 -10564 -1018 -10530
rect -860 -10564 -826 -10530
rect -668 -10564 -634 -10530
rect -476 -10564 -442 -10530
rect -284 -10564 -250 -10530
rect -92 -10564 -58 -10530
rect 100 -10564 134 -10530
rect 292 -10564 326 -10530
rect 484 -10564 518 -10530
rect 676 -10564 710 -10530
rect 868 -10564 902 -10530
rect 1060 -10564 1094 -10530
rect -1052 -10672 -1018 -10638
rect -860 -10672 -826 -10638
rect -668 -10672 -634 -10638
rect -476 -10672 -442 -10638
rect -284 -10672 -250 -10638
rect -92 -10672 -58 -10638
rect 100 -10672 134 -10638
rect 292 -10672 326 -10638
rect 484 -10672 518 -10638
rect 676 -10672 710 -10638
rect 868 -10672 902 -10638
rect 1060 -10672 1094 -10638
rect -1148 -11182 -1114 -11148
rect -956 -11182 -922 -11148
rect -764 -11182 -730 -11148
rect -572 -11182 -538 -11148
rect -380 -11182 -346 -11148
rect -188 -11182 -154 -11148
rect 4 -11182 38 -11148
rect 196 -11182 230 -11148
rect 388 -11182 422 -11148
rect 580 -11182 614 -11148
rect 772 -11182 806 -11148
rect 964 -11182 998 -11148
rect 1156 -11182 1190 -11148
rect 1676 -8872 1844 -8838
rect 1934 -8872 2102 -8838
rect 2192 -8872 2360 -8838
rect 2450 -8872 2618 -8838
rect 2708 -8872 2876 -8838
rect 2966 -8872 3134 -8838
rect 1676 -9382 1844 -9348
rect 1934 -9382 2102 -9348
rect 2192 -9382 2360 -9348
rect 2450 -9382 2618 -9348
rect 2708 -9382 2876 -9348
rect 2966 -9382 3134 -9348
rect 3572 -8872 3740 -8838
rect 3830 -8872 3998 -8838
rect 4088 -8872 4256 -8838
rect 4346 -8872 4514 -8838
rect 4604 -8872 4772 -8838
rect 4862 -8872 5030 -8838
rect 3572 -9382 3740 -9348
rect 3830 -9382 3998 -9348
rect 4088 -9382 4256 -9348
rect 4346 -9382 4514 -9348
rect 4604 -9382 4772 -9348
rect 4862 -9382 5030 -9348
rect 5604 -8872 5638 -8838
rect 5796 -8872 5830 -8838
rect 5508 -9382 5542 -9348
rect 5700 -9382 5734 -9348
rect 5892 -9382 5926 -9348
rect 1709 -9884 2077 -9850
rect 2629 -9884 2997 -9850
rect 3549 -9884 3917 -9850
rect 4469 -9884 4837 -9850
rect 5389 -9884 5757 -9850
rect 1709 -10994 2077 -10960
rect 2629 -10994 2997 -10960
rect 3549 -10994 3917 -10960
rect 4469 -10994 4837 -10960
rect 5389 -10994 5757 -10960
rect 6392 -10164 6560 -10130
rect 6392 -10392 6560 -10358
rect 6392 -10732 6560 -10698
rect 6392 -10942 6560 -10908
<< locali >>
rect -1296 2728 2324 2790
rect -1296 2710 -1194 2728
rect -1290 2694 -1194 2710
rect 346 2694 604 2728
rect 2144 2694 2324 2728
rect -1290 2632 -1256 2694
rect 408 2632 542 2694
rect -1143 2592 -1127 2626
rect -1093 2592 -1029 2626
rect -995 2592 -931 2626
rect -897 2592 -833 2626
rect -799 2592 -735 2626
rect -701 2592 -637 2626
rect -603 2592 -539 2626
rect -505 2592 -441 2626
rect -407 2592 -343 2626
rect -309 2592 -245 2626
rect -211 2592 -147 2626
rect -113 2592 -49 2626
rect -15 2592 49 2626
rect 83 2592 147 2626
rect 181 2592 245 2626
rect 279 2592 295 2626
rect -1176 2533 -1142 2549
rect -1176 2141 -1142 2157
rect -1078 2533 -1044 2549
rect -1078 2141 -1044 2157
rect -980 2533 -946 2549
rect -980 2141 -946 2157
rect -882 2533 -848 2549
rect -882 2141 -848 2157
rect -784 2533 -750 2549
rect -784 2141 -750 2157
rect -686 2533 -652 2549
rect -686 2141 -652 2157
rect -588 2533 -554 2549
rect -588 2141 -554 2157
rect -490 2533 -456 2549
rect -490 2141 -456 2157
rect -392 2533 -358 2549
rect -392 2141 -358 2157
rect -294 2533 -260 2549
rect -294 2141 -260 2157
rect -196 2533 -162 2549
rect -196 2141 -162 2157
rect -98 2533 -64 2549
rect -98 2141 -64 2157
rect 0 2533 34 2549
rect 0 2141 34 2157
rect 98 2533 132 2549
rect 98 2141 132 2157
rect 196 2533 230 2549
rect 196 2141 230 2157
rect 294 2533 328 2549
rect 294 2141 328 2157
rect -1143 2064 -1127 2098
rect -1093 2064 -1029 2098
rect -995 2064 -931 2098
rect -897 2064 -833 2098
rect -799 2064 -735 2098
rect -701 2064 -637 2098
rect -603 2064 -539 2098
rect -505 2064 -441 2098
rect -407 2064 -343 2098
rect -309 2064 -245 2098
rect -211 2064 -147 2098
rect -113 2064 -49 2098
rect -15 2064 49 2098
rect 83 2064 147 2098
rect 181 2064 245 2098
rect 279 2064 295 2098
rect -1143 1956 -1127 1990
rect -1093 1956 -1029 1990
rect -995 1956 -931 1990
rect -897 1956 -833 1990
rect -799 1956 -735 1990
rect -701 1956 -637 1990
rect -603 1956 -539 1990
rect -505 1956 -441 1990
rect -407 1956 -343 1990
rect -309 1956 -245 1990
rect -211 1956 -147 1990
rect -113 1956 -49 1990
rect -15 1956 49 1990
rect 83 1956 147 1990
rect 181 1956 245 1990
rect 279 1956 295 1990
rect -1176 1897 -1142 1913
rect -1176 1505 -1142 1521
rect -1078 1897 -1044 1913
rect -1078 1505 -1044 1521
rect -980 1897 -946 1913
rect -980 1505 -946 1521
rect -882 1897 -848 1913
rect -882 1505 -848 1521
rect -784 1897 -750 1913
rect -784 1505 -750 1521
rect -686 1897 -652 1913
rect -686 1505 -652 1521
rect -588 1897 -554 1913
rect -588 1505 -554 1521
rect -490 1897 -456 1913
rect -490 1505 -456 1521
rect -392 1897 -358 1913
rect -392 1505 -358 1521
rect -294 1897 -260 1913
rect -294 1505 -260 1521
rect -196 1897 -162 1913
rect -196 1505 -162 1521
rect -98 1897 -64 1913
rect -98 1505 -64 1521
rect 0 1897 34 1913
rect 0 1505 34 1521
rect 98 1897 132 1913
rect 98 1505 132 1521
rect 196 1897 230 1913
rect 196 1505 230 1521
rect 294 1897 328 1913
rect 294 1505 328 1521
rect -1143 1428 -1127 1462
rect -1093 1428 -1029 1462
rect -995 1428 -931 1462
rect -897 1428 -833 1462
rect -799 1428 -735 1462
rect -701 1428 -637 1462
rect -603 1428 -539 1462
rect -505 1428 -441 1462
rect -407 1428 -343 1462
rect -309 1428 -245 1462
rect -211 1428 -147 1462
rect -113 1428 -49 1462
rect -15 1428 49 1462
rect 83 1428 147 1462
rect 181 1428 245 1462
rect 279 1428 295 1462
rect -1290 1360 -1256 1422
rect 442 1422 508 2632
rect 2206 2632 2324 2694
rect 655 2592 671 2626
rect 705 2592 769 2626
rect 803 2592 867 2626
rect 901 2592 965 2626
rect 999 2592 1063 2626
rect 1097 2592 1161 2626
rect 1195 2592 1259 2626
rect 1293 2592 1357 2626
rect 1391 2592 1455 2626
rect 1489 2592 1553 2626
rect 1587 2592 1651 2626
rect 1685 2592 1749 2626
rect 1783 2592 1847 2626
rect 1881 2592 1945 2626
rect 1979 2592 2043 2626
rect 2077 2592 2093 2626
rect 622 2533 656 2549
rect 622 2141 656 2157
rect 720 2533 754 2549
rect 720 2141 754 2157
rect 818 2533 852 2549
rect 818 2141 852 2157
rect 916 2533 950 2549
rect 916 2141 950 2157
rect 1014 2533 1048 2549
rect 1014 2141 1048 2157
rect 1112 2533 1146 2549
rect 1112 2141 1146 2157
rect 1210 2533 1244 2549
rect 1210 2141 1244 2157
rect 1308 2533 1342 2549
rect 1308 2141 1342 2157
rect 1406 2533 1440 2549
rect 1406 2141 1440 2157
rect 1504 2533 1538 2549
rect 1504 2141 1538 2157
rect 1602 2533 1636 2549
rect 1602 2141 1636 2157
rect 1700 2533 1734 2549
rect 1700 2141 1734 2157
rect 1798 2533 1832 2549
rect 1798 2141 1832 2157
rect 1896 2533 1930 2549
rect 1896 2141 1930 2157
rect 1994 2533 2028 2549
rect 1994 2141 2028 2157
rect 2092 2533 2126 2549
rect 2092 2141 2126 2157
rect 655 2064 671 2098
rect 705 2064 769 2098
rect 803 2064 867 2098
rect 901 2064 965 2098
rect 999 2064 1063 2098
rect 1097 2064 1161 2098
rect 1195 2064 1259 2098
rect 1293 2064 1357 2098
rect 1391 2064 1455 2098
rect 1489 2064 1553 2098
rect 1587 2064 1651 2098
rect 1685 2064 1749 2098
rect 1783 2064 1847 2098
rect 1881 2064 1945 2098
rect 1979 2064 2043 2098
rect 2077 2064 2093 2098
rect 2240 2160 2324 2632
rect 2240 2076 4394 2160
rect 2240 2070 2406 2076
rect 655 1956 671 1990
rect 705 1956 769 1990
rect 803 1956 867 1990
rect 901 1956 965 1990
rect 999 1956 1063 1990
rect 1097 1956 1161 1990
rect 1195 1956 1259 1990
rect 1293 1956 1357 1990
rect 1391 1956 1455 1990
rect 1489 1956 1553 1990
rect 1587 1956 1651 1990
rect 1685 1956 1749 1990
rect 1783 1956 1847 1990
rect 1881 1956 1945 1990
rect 1979 1956 2043 1990
rect 2077 1956 2093 1990
rect 622 1897 656 1913
rect 622 1505 656 1521
rect 720 1897 754 1913
rect 720 1505 754 1521
rect 818 1897 852 1913
rect 818 1505 852 1521
rect 916 1897 950 1913
rect 916 1505 950 1521
rect 1014 1897 1048 1913
rect 1014 1505 1048 1521
rect 1112 1897 1146 1913
rect 1112 1505 1146 1521
rect 1210 1897 1244 1913
rect 1210 1505 1244 1521
rect 1308 1897 1342 1913
rect 1308 1505 1342 1521
rect 1406 1897 1440 1913
rect 1406 1505 1440 1521
rect 1504 1897 1538 1913
rect 1504 1505 1538 1521
rect 1602 1897 1636 1913
rect 1602 1505 1636 1521
rect 1700 1897 1734 1913
rect 1700 1505 1734 1521
rect 1798 1897 1832 1913
rect 1798 1505 1832 1521
rect 1896 1897 1930 1913
rect 1896 1505 1930 1521
rect 1994 1897 2028 1913
rect 1994 1505 2028 1521
rect 2092 1897 2126 1913
rect 2092 1505 2126 1521
rect 2344 2042 2406 2070
rect 4056 2042 4394 2076
rect 4118 1980 4394 2042
rect 2470 1940 2486 1974
rect 2554 1940 2570 1974
rect 2628 1940 2644 1974
rect 2712 1940 2728 1974
rect 2786 1940 2802 1974
rect 2870 1940 2886 1974
rect 2944 1940 2960 1974
rect 3028 1940 3044 1974
rect 3102 1940 3118 1974
rect 3186 1940 3202 1974
rect 3260 1940 3276 1974
rect 3344 1940 3360 1974
rect 3418 1940 3434 1974
rect 3502 1940 3518 1974
rect 3576 1940 3592 1974
rect 3660 1940 3676 1974
rect 3734 1940 3750 1974
rect 3818 1940 3834 1974
rect 3892 1940 3908 1974
rect 3976 1940 3992 1974
rect 655 1428 671 1462
rect 705 1428 769 1462
rect 803 1428 867 1462
rect 901 1428 965 1462
rect 999 1428 1063 1462
rect 1097 1428 1161 1462
rect 1195 1428 1259 1462
rect 1293 1428 1357 1462
rect 1391 1428 1455 1462
rect 1489 1428 1553 1462
rect 1587 1428 1651 1462
rect 1685 1428 1749 1462
rect 1783 1428 1847 1462
rect 1881 1428 1945 1462
rect 1979 1428 2043 1462
rect 2077 1428 2093 1462
rect 408 1360 542 1422
rect 2240 1422 2310 1510
rect 2206 1406 2310 1422
rect 2424 1881 2458 1897
rect 2424 1489 2458 1505
rect 2582 1881 2616 1897
rect 2582 1489 2616 1505
rect 2740 1881 2774 1897
rect 2740 1489 2774 1505
rect 2898 1881 2932 1897
rect 2898 1489 2932 1505
rect 3056 1881 3090 1897
rect 3056 1489 3090 1505
rect 3214 1881 3248 1897
rect 3214 1489 3248 1505
rect 3372 1881 3406 1897
rect 3372 1489 3406 1505
rect 3530 1881 3564 1897
rect 3530 1489 3564 1505
rect 3688 1881 3722 1897
rect 3688 1489 3722 1505
rect 3846 1881 3880 1897
rect 3846 1489 3880 1505
rect 4004 1881 4038 1897
rect 4004 1489 4038 1505
rect 2470 1412 2486 1446
rect 2554 1412 2570 1446
rect 2628 1412 2644 1446
rect 2712 1412 2728 1446
rect 2786 1412 2802 1446
rect 2870 1412 2886 1446
rect 2944 1412 2960 1446
rect 3028 1412 3044 1446
rect 3102 1412 3118 1446
rect 3186 1412 3202 1446
rect 3260 1412 3276 1446
rect 3344 1412 3360 1446
rect 3418 1412 3434 1446
rect 3502 1412 3518 1446
rect 3576 1412 3592 1446
rect 3660 1412 3676 1446
rect 3734 1412 3750 1446
rect 3818 1412 3834 1446
rect 3892 1412 3908 1446
rect 3976 1412 3992 1446
rect 2206 1360 2344 1406
rect -1290 1326 -1194 1360
rect 346 1330 604 1360
rect 346 1326 442 1330
rect 508 1326 604 1330
rect 2144 1344 2344 1360
rect 4152 1406 4394 1980
rect 4118 1344 4394 1406
rect 2144 1326 2406 1344
rect 2074 1310 2406 1326
rect 4056 1310 4394 1344
rect -1290 1240 -1194 1252
rect -1396 1218 -1194 1240
rect 1326 1250 1422 1252
rect 1326 1218 1534 1250
rect 2074 1233 4394 1310
rect -1396 1156 -1256 1218
rect -1396 -18 -1290 1156
rect 1388 1156 1534 1218
rect -1144 1116 -1127 1150
rect -1093 1116 -1030 1150
rect -996 1116 -931 1150
rect -897 1116 -834 1150
rect -800 1116 -735 1150
rect -701 1116 -638 1150
rect -604 1116 -539 1150
rect -505 1116 -442 1150
rect -408 1116 -343 1150
rect -309 1116 -246 1150
rect -212 1116 -147 1150
rect -113 1116 -50 1150
rect -16 1116 49 1150
rect 83 1116 146 1150
rect 180 1116 245 1150
rect 279 1116 342 1150
rect 376 1116 441 1150
rect 475 1116 538 1150
rect 572 1116 637 1150
rect 671 1116 734 1150
rect 768 1116 833 1150
rect 867 1116 930 1150
rect 964 1116 1029 1150
rect 1063 1116 1126 1150
rect 1160 1116 1225 1150
rect 1259 1116 1275 1150
rect -1176 1066 -1142 1082
rect -1176 674 -1142 690
rect -1078 1066 -1044 1082
rect -1078 674 -1044 690
rect -980 1066 -946 1082
rect -980 674 -946 690
rect -882 1066 -848 1082
rect -882 674 -848 690
rect -784 1066 -750 1082
rect -784 674 -750 690
rect -686 1066 -652 1082
rect -686 674 -652 690
rect -588 1066 -554 1082
rect -588 674 -554 690
rect -490 1066 -456 1082
rect -490 674 -456 690
rect -392 1066 -358 1082
rect -392 674 -358 690
rect -294 1066 -260 1082
rect -294 674 -260 690
rect -196 1066 -162 1082
rect -196 674 -162 690
rect -98 1066 -64 1082
rect -98 674 -64 690
rect 0 1066 34 1082
rect 0 674 34 690
rect 98 1066 132 1082
rect 98 674 132 690
rect 196 1066 230 1082
rect 196 674 230 690
rect 294 1066 328 1082
rect 294 674 328 690
rect 392 1066 426 1082
rect 392 674 426 690
rect 490 1066 524 1082
rect 490 674 524 690
rect 588 1066 622 1082
rect 588 674 622 690
rect 686 1066 720 1082
rect 686 674 720 690
rect 784 1066 818 1082
rect 784 674 818 690
rect 882 1066 916 1082
rect 882 674 916 690
rect 980 1066 1014 1082
rect 980 674 1014 690
rect 1078 1066 1112 1082
rect 1078 674 1112 690
rect 1176 1066 1210 1082
rect 1176 674 1210 690
rect 1274 1066 1308 1082
rect 1274 674 1308 690
rect -1144 606 -1128 640
rect -1094 606 -1029 640
rect -995 606 -932 640
rect -898 606 -833 640
rect -799 606 -736 640
rect -702 606 -637 640
rect -603 606 -540 640
rect -506 606 -441 640
rect -407 606 -344 640
rect -310 606 -245 640
rect -211 606 -148 640
rect -114 606 -49 640
rect -15 606 48 640
rect 82 606 147 640
rect 181 606 244 640
rect 278 606 343 640
rect 377 606 440 640
rect 474 606 539 640
rect 573 606 636 640
rect 670 606 735 640
rect 769 606 832 640
rect 866 606 931 640
rect 965 606 1028 640
rect 1062 606 1127 640
rect 1161 606 1224 640
rect 1258 606 1274 640
rect -1143 498 -1127 532
rect -1093 498 -1029 532
rect -995 498 -931 532
rect -897 498 -833 532
rect -799 498 -735 532
rect -701 498 -637 532
rect -603 498 -539 532
rect -505 498 -441 532
rect -407 498 -343 532
rect -309 498 -245 532
rect -211 498 -147 532
rect -113 498 -49 532
rect -15 498 49 532
rect 83 498 147 532
rect 181 498 245 532
rect 279 498 343 532
rect 377 498 441 532
rect 475 498 539 532
rect 573 498 637 532
rect 671 498 735 532
rect 769 498 833 532
rect 867 498 931 532
rect 965 498 1029 532
rect 1063 498 1127 532
rect 1161 498 1225 532
rect 1259 498 1275 532
rect -1176 448 -1142 464
rect -1176 56 -1142 72
rect -1078 448 -1044 464
rect -1078 56 -1044 72
rect -980 448 -946 464
rect -980 56 -946 72
rect -882 448 -848 464
rect -882 56 -848 72
rect -784 448 -750 464
rect -784 56 -750 72
rect -686 448 -652 464
rect -686 56 -652 72
rect -588 448 -554 464
rect -588 56 -554 72
rect -490 448 -456 464
rect -490 56 -456 72
rect -392 448 -358 464
rect -392 56 -358 72
rect -294 448 -260 464
rect -294 56 -260 72
rect -196 448 -162 464
rect -196 56 -162 72
rect -98 448 -64 464
rect -98 56 -64 72
rect 0 448 34 464
rect 0 56 34 72
rect 98 448 132 464
rect 98 56 132 72
rect 196 448 230 464
rect 196 56 230 72
rect 294 448 328 464
rect 294 56 328 72
rect 392 448 426 464
rect 392 56 426 72
rect 490 448 524 464
rect 490 56 524 72
rect 588 448 622 464
rect 588 56 622 72
rect 686 448 720 464
rect 686 56 720 72
rect 784 448 818 464
rect 784 56 818 72
rect 882 448 916 464
rect 882 56 916 72
rect 980 448 1014 464
rect 980 56 1014 72
rect 1078 448 1112 464
rect 1078 56 1112 72
rect 1176 448 1210 464
rect 1176 56 1210 72
rect 1274 448 1308 464
rect 1274 56 1308 72
rect -1143 -12 -1127 22
rect -1093 -12 -1029 22
rect -995 -12 -931 22
rect -897 -12 -833 22
rect -799 -12 -735 22
rect -701 -12 -637 22
rect -603 -12 -539 22
rect -505 -12 -441 22
rect -407 -12 -343 22
rect -309 -12 -245 22
rect -211 -12 -147 22
rect -113 -12 -49 22
rect -15 -12 49 22
rect 83 -12 147 22
rect 181 -12 245 22
rect 279 -12 343 22
rect 377 -12 441 22
rect 475 -12 539 22
rect 573 -12 637 22
rect 671 -12 735 22
rect 769 -12 833 22
rect 867 -12 931 22
rect 965 -12 1029 22
rect 1063 -12 1127 22
rect 1161 -12 1225 22
rect 1259 -12 1275 22
rect -1396 -80 -1256 -18
rect 1422 -18 1534 1156
rect 1388 -80 1534 -18
rect -1396 -114 -1194 -80
rect 1326 -114 1534 -80
rect -1396 -192 1534 -114
rect -1396 -226 -1194 -192
rect 1326 -226 1534 -192
rect -1396 -288 -1256 -226
rect -1396 -1462 -1290 -288
rect 1388 -288 1534 -226
rect -1144 -328 -1127 -294
rect -1093 -328 -1030 -294
rect -996 -328 -931 -294
rect -897 -328 -834 -294
rect -800 -328 -735 -294
rect -701 -328 -638 -294
rect -604 -328 -539 -294
rect -505 -328 -442 -294
rect -408 -328 -343 -294
rect -309 -328 -246 -294
rect -212 -328 -147 -294
rect -113 -328 -50 -294
rect -16 -328 49 -294
rect 83 -328 146 -294
rect 180 -328 245 -294
rect 279 -328 342 -294
rect 376 -328 441 -294
rect 475 -328 538 -294
rect 572 -328 637 -294
rect 671 -328 734 -294
rect 768 -328 833 -294
rect 867 -328 930 -294
rect 964 -328 1029 -294
rect 1063 -328 1126 -294
rect 1160 -328 1225 -294
rect 1259 -328 1275 -294
rect -1176 -378 -1142 -362
rect -1176 -770 -1142 -754
rect -1078 -378 -1044 -362
rect -1078 -770 -1044 -754
rect -980 -378 -946 -362
rect -980 -770 -946 -754
rect -882 -378 -848 -362
rect -882 -770 -848 -754
rect -784 -378 -750 -362
rect -784 -770 -750 -754
rect -686 -378 -652 -362
rect -686 -770 -652 -754
rect -588 -378 -554 -362
rect -588 -770 -554 -754
rect -490 -378 -456 -362
rect -490 -770 -456 -754
rect -392 -378 -358 -362
rect -392 -770 -358 -754
rect -294 -378 -260 -362
rect -294 -770 -260 -754
rect -196 -378 -162 -362
rect -196 -770 -162 -754
rect -98 -378 -64 -362
rect -98 -770 -64 -754
rect 0 -378 34 -362
rect 0 -770 34 -754
rect 98 -378 132 -362
rect 98 -770 132 -754
rect 196 -378 230 -362
rect 196 -770 230 -754
rect 294 -378 328 -362
rect 294 -770 328 -754
rect 392 -378 426 -362
rect 392 -770 426 -754
rect 490 -378 524 -362
rect 490 -770 524 -754
rect 588 -378 622 -362
rect 588 -770 622 -754
rect 686 -378 720 -362
rect 686 -770 720 -754
rect 784 -378 818 -362
rect 784 -770 818 -754
rect 882 -378 916 -362
rect 882 -770 916 -754
rect 980 -378 1014 -362
rect 980 -770 1014 -754
rect 1078 -378 1112 -362
rect 1078 -770 1112 -754
rect 1176 -378 1210 -362
rect 1176 -770 1210 -754
rect 1274 -378 1308 -362
rect 1274 -770 1308 -754
rect -1144 -838 -1128 -804
rect -1094 -838 -1029 -804
rect -995 -838 -932 -804
rect -898 -838 -833 -804
rect -799 -838 -736 -804
rect -702 -838 -637 -804
rect -603 -838 -540 -804
rect -506 -838 -441 -804
rect -407 -838 -344 -804
rect -310 -838 -245 -804
rect -211 -838 -148 -804
rect -114 -838 -49 -804
rect -15 -838 48 -804
rect 82 -838 147 -804
rect 181 -838 244 -804
rect 278 -838 343 -804
rect 377 -838 440 -804
rect 474 -838 539 -804
rect 573 -838 636 -804
rect 670 -838 735 -804
rect 769 -838 832 -804
rect 866 -838 931 -804
rect 965 -838 1028 -804
rect 1062 -838 1127 -804
rect 1161 -838 1224 -804
rect 1258 -838 1274 -804
rect -1143 -946 -1127 -912
rect -1093 -946 -1029 -912
rect -995 -946 -931 -912
rect -897 -946 -833 -912
rect -799 -946 -735 -912
rect -701 -946 -637 -912
rect -603 -946 -539 -912
rect -505 -946 -441 -912
rect -407 -946 -343 -912
rect -309 -946 -245 -912
rect -211 -946 -147 -912
rect -113 -946 -49 -912
rect -15 -946 49 -912
rect 83 -946 147 -912
rect 181 -946 245 -912
rect 279 -946 343 -912
rect 377 -946 441 -912
rect 475 -946 539 -912
rect 573 -946 637 -912
rect 671 -946 735 -912
rect 769 -946 833 -912
rect 867 -946 931 -912
rect 965 -946 1029 -912
rect 1063 -946 1127 -912
rect 1161 -946 1225 -912
rect 1259 -946 1275 -912
rect -1176 -996 -1142 -980
rect -1176 -1388 -1142 -1372
rect -1078 -996 -1044 -980
rect -1078 -1388 -1044 -1372
rect -980 -996 -946 -980
rect -980 -1388 -946 -1372
rect -882 -996 -848 -980
rect -882 -1388 -848 -1372
rect -784 -996 -750 -980
rect -784 -1388 -750 -1372
rect -686 -996 -652 -980
rect -686 -1388 -652 -1372
rect -588 -996 -554 -980
rect -588 -1388 -554 -1372
rect -490 -996 -456 -980
rect -490 -1388 -456 -1372
rect -392 -996 -358 -980
rect -392 -1388 -358 -1372
rect -294 -996 -260 -980
rect -294 -1388 -260 -1372
rect -196 -996 -162 -980
rect -196 -1388 -162 -1372
rect -98 -996 -64 -980
rect -98 -1388 -64 -1372
rect 0 -996 34 -980
rect 0 -1388 34 -1372
rect 98 -996 132 -980
rect 98 -1388 132 -1372
rect 196 -996 230 -980
rect 196 -1388 230 -1372
rect 294 -996 328 -980
rect 294 -1388 328 -1372
rect 392 -996 426 -980
rect 392 -1388 426 -1372
rect 490 -996 524 -980
rect 490 -1388 524 -1372
rect 588 -996 622 -980
rect 588 -1388 622 -1372
rect 686 -996 720 -980
rect 686 -1388 720 -1372
rect 784 -996 818 -980
rect 784 -1388 818 -1372
rect 882 -996 916 -980
rect 882 -1388 916 -1372
rect 980 -996 1014 -980
rect 980 -1388 1014 -1372
rect 1078 -996 1112 -980
rect 1078 -1388 1112 -1372
rect 1176 -996 1210 -980
rect 1176 -1388 1210 -1372
rect 1274 -996 1308 -980
rect 1274 -1388 1308 -1372
rect -1143 -1456 -1127 -1422
rect -1093 -1456 -1029 -1422
rect -995 -1456 -931 -1422
rect -897 -1456 -833 -1422
rect -799 -1456 -735 -1422
rect -701 -1456 -637 -1422
rect -603 -1456 -539 -1422
rect -505 -1456 -441 -1422
rect -407 -1456 -343 -1422
rect -309 -1456 -245 -1422
rect -211 -1456 -147 -1422
rect -113 -1456 -49 -1422
rect -15 -1456 49 -1422
rect 83 -1456 147 -1422
rect 181 -1456 245 -1422
rect 279 -1456 343 -1422
rect 377 -1456 441 -1422
rect 475 -1456 539 -1422
rect 573 -1456 637 -1422
rect 671 -1456 735 -1422
rect 769 -1456 833 -1422
rect 867 -1456 931 -1422
rect 965 -1456 1029 -1422
rect 1063 -1456 1127 -1422
rect 1161 -1456 1225 -1422
rect 1259 -1456 1275 -1422
rect -1396 -1524 -1256 -1462
rect 1422 -846 1534 -288
rect 2071 1199 2131 1233
rect 4337 1199 4397 1233
rect 2071 1173 2105 1199
rect 4363 1173 4397 1199
rect 2304 932 4174 1000
rect 2304 898 2466 932
rect 4006 898 4174 932
rect 2304 836 2404 898
rect 2304 320 2370 836
rect 2284 160 2370 320
rect 2294 -338 2370 160
rect 4068 836 4174 898
rect 2517 796 2533 830
rect 2567 796 2631 830
rect 2665 796 2729 830
rect 2763 796 2827 830
rect 2861 796 2925 830
rect 2959 796 3023 830
rect 3057 796 3121 830
rect 3155 796 3219 830
rect 3253 796 3317 830
rect 3351 796 3415 830
rect 3449 796 3513 830
rect 3547 796 3611 830
rect 3645 796 3709 830
rect 3743 796 3807 830
rect 3841 796 3905 830
rect 3939 796 3955 830
rect 2484 746 2518 762
rect 2484 354 2518 370
rect 2582 746 2616 762
rect 2582 354 2616 370
rect 2680 746 2714 762
rect 2680 354 2714 370
rect 2778 746 2812 762
rect 2778 354 2812 370
rect 2876 746 2910 762
rect 2876 354 2910 370
rect 2974 746 3008 762
rect 2974 354 3008 370
rect 3072 746 3106 762
rect 3072 354 3106 370
rect 3170 746 3204 762
rect 3170 354 3204 370
rect 3268 746 3302 762
rect 3268 354 3302 370
rect 3366 746 3400 762
rect 3366 354 3400 370
rect 3464 746 3498 762
rect 3464 354 3498 370
rect 3562 746 3596 762
rect 3562 354 3596 370
rect 3660 746 3694 762
rect 3660 354 3694 370
rect 3758 746 3792 762
rect 3758 354 3792 370
rect 3856 746 3890 762
rect 3856 354 3890 370
rect 3954 746 3988 762
rect 3954 354 3988 370
rect 4102 340 4174 836
rect 2517 286 2533 320
rect 2567 286 2631 320
rect 2665 286 2729 320
rect 2763 286 2827 320
rect 2861 286 2925 320
rect 2959 286 3023 320
rect 3057 286 3121 320
rect 3155 286 3219 320
rect 3253 286 3317 320
rect 3351 286 3415 320
rect 3449 286 3513 320
rect 3547 286 3611 320
rect 3645 286 3709 320
rect 3743 286 3807 320
rect 3841 286 3905 320
rect 3939 286 3955 320
rect 2517 178 2533 212
rect 2567 178 2631 212
rect 2665 178 2729 212
rect 2763 178 2827 212
rect 2861 178 2925 212
rect 2959 178 3023 212
rect 3057 178 3121 212
rect 3155 178 3219 212
rect 3253 178 3317 212
rect 3351 178 3415 212
rect 3449 178 3513 212
rect 3547 178 3611 212
rect 3645 178 3709 212
rect 3743 178 3807 212
rect 3841 178 3905 212
rect 3939 178 3955 212
rect 2484 128 2518 144
rect 2484 -264 2518 -248
rect 2582 128 2616 144
rect 2582 -264 2616 -248
rect 2680 128 2714 144
rect 2680 -264 2714 -248
rect 2778 128 2812 144
rect 2778 -264 2812 -248
rect 2876 128 2910 144
rect 2876 -264 2910 -248
rect 2974 128 3008 144
rect 2974 -264 3008 -248
rect 3072 128 3106 144
rect 3072 -264 3106 -248
rect 3170 128 3204 144
rect 3170 -264 3204 -248
rect 3268 128 3302 144
rect 3268 -264 3302 -248
rect 3366 128 3400 144
rect 3366 -264 3400 -248
rect 3464 128 3498 144
rect 3464 -264 3498 -248
rect 3562 128 3596 144
rect 3562 -264 3596 -248
rect 3660 128 3694 144
rect 3660 -264 3694 -248
rect 3758 128 3792 144
rect 3758 -264 3792 -248
rect 3856 128 3890 144
rect 3856 -264 3890 -248
rect 3954 128 3988 144
rect 3954 -264 3988 -248
rect 2517 -332 2533 -298
rect 2567 -332 2631 -298
rect 2665 -332 2729 -298
rect 2763 -332 2827 -298
rect 2861 -332 2925 -298
rect 2959 -332 3023 -298
rect 3057 -332 3121 -298
rect 3155 -332 3219 -298
rect 3253 -332 3317 -298
rect 3351 -332 3415 -298
rect 3449 -332 3513 -298
rect 3547 -332 3611 -298
rect 3645 -332 3709 -298
rect 3743 -332 3807 -298
rect 3841 -332 3905 -298
rect 3939 -332 3955 -298
rect 2294 -400 2404 -338
rect 4102 -338 4174 130
rect 4068 -400 4174 -338
rect 2294 -434 2466 -400
rect 4006 -434 4174 -400
rect 2294 -500 4174 -434
rect 2071 -699 2105 -673
rect 4363 -699 4397 -673
rect 2071 -733 2131 -699
rect 4337 -733 4397 -699
rect 1422 -880 1596 -846
rect 2818 -880 2914 -846
rect 1422 -942 1534 -880
rect 1422 -1462 1500 -942
rect 1388 -1498 1500 -1462
rect 2880 -942 2914 -880
rect 1646 -982 1662 -948
rect 1696 -982 1758 -948
rect 1792 -982 1854 -948
rect 1888 -982 1950 -948
rect 1984 -982 2046 -948
rect 2080 -982 2142 -948
rect 2176 -982 2238 -948
rect 2272 -982 2334 -948
rect 2368 -982 2430 -948
rect 2464 -982 2526 -948
rect 2560 -982 2622 -948
rect 2656 -982 2718 -948
rect 2752 -982 2768 -948
rect 1614 -1032 1648 -1016
rect 1614 -1424 1648 -1408
rect 1710 -1032 1744 -1016
rect 1710 -1424 1744 -1408
rect 1806 -1032 1840 -1016
rect 1806 -1424 1840 -1408
rect 1902 -1032 1936 -1016
rect 1902 -1424 1936 -1408
rect 1998 -1032 2032 -1016
rect 1998 -1424 2032 -1408
rect 2094 -1032 2128 -1016
rect 2094 -1424 2128 -1408
rect 2190 -1032 2224 -1016
rect 2190 -1424 2224 -1408
rect 2286 -1032 2320 -1016
rect 2286 -1424 2320 -1408
rect 2382 -1032 2416 -1016
rect 2382 -1424 2416 -1408
rect 2478 -1032 2512 -1016
rect 2478 -1424 2512 -1408
rect 2574 -1032 2608 -1016
rect 2574 -1424 2608 -1408
rect 2670 -1032 2704 -1016
rect 2670 -1424 2704 -1408
rect 2766 -1032 2800 -1016
rect 2766 -1424 2800 -1408
rect 1646 -1492 1662 -1458
rect 1696 -1492 1758 -1458
rect 1792 -1492 1854 -1458
rect 1888 -1492 1950 -1458
rect 1984 -1492 2046 -1458
rect 2080 -1492 2142 -1458
rect 2176 -1492 2238 -1458
rect 2272 -1492 2334 -1458
rect 2368 -1492 2430 -1458
rect 2464 -1492 2526 -1458
rect 2560 -1492 2622 -1458
rect 2656 -1492 2718 -1458
rect 2752 -1492 2768 -1458
rect 1388 -1524 1534 -1498
rect -1396 -1558 -1194 -1524
rect 1326 -1558 1534 -1524
rect -1396 -1560 1534 -1558
rect 2880 -1560 2914 -1498
rect -1396 -1594 1596 -1560
rect 2818 -1594 2914 -1560
rect -1396 -1612 2914 -1594
rect -1396 -1646 -1214 -1612
rect 1256 -1646 2914 -1612
rect -1396 -1708 -1256 -1646
rect -1396 -4118 -1310 -1708
rect -1276 -4118 -1256 -1708
rect 1318 -1666 2914 -1646
rect 1318 -1700 1596 -1666
rect 3214 -1700 3310 -1666
rect 1318 -1708 1534 -1700
rect -1164 -1748 -1148 -1714
rect -1114 -1748 -1098 -1714
rect -972 -1748 -956 -1714
rect -922 -1748 -906 -1714
rect -780 -1748 -764 -1714
rect -730 -1748 -714 -1714
rect -588 -1748 -572 -1714
rect -538 -1748 -522 -1714
rect -396 -1748 -380 -1714
rect -346 -1748 -330 -1714
rect -204 -1748 -188 -1714
rect -154 -1748 -138 -1714
rect -12 -1748 4 -1714
rect 38 -1748 54 -1714
rect 180 -1748 196 -1714
rect 230 -1748 246 -1714
rect 372 -1748 388 -1714
rect 422 -1748 438 -1714
rect 564 -1748 580 -1714
rect 614 -1748 630 -1714
rect 756 -1748 772 -1714
rect 806 -1748 822 -1714
rect 948 -1748 964 -1714
rect 998 -1748 1014 -1714
rect 1140 -1748 1156 -1714
rect 1190 -1748 1206 -1714
rect -1196 -1798 -1162 -1782
rect -1196 -2190 -1162 -2174
rect -1100 -1798 -1066 -1782
rect -1100 -2190 -1066 -2174
rect -1004 -1798 -970 -1782
rect -1004 -2190 -970 -2174
rect -908 -1798 -874 -1782
rect -908 -2190 -874 -2174
rect -812 -1798 -778 -1782
rect -812 -2190 -778 -2174
rect -716 -1798 -682 -1782
rect -716 -2190 -682 -2174
rect -620 -1798 -586 -1782
rect -620 -2190 -586 -2174
rect -524 -1798 -490 -1782
rect -524 -2190 -490 -2174
rect -428 -1798 -394 -1782
rect -428 -2190 -394 -2174
rect -332 -1798 -298 -1782
rect -332 -2190 -298 -2174
rect -236 -1798 -202 -1782
rect -236 -2190 -202 -2174
rect -140 -1798 -106 -1782
rect -140 -2190 -106 -2174
rect -44 -1798 -10 -1782
rect -44 -2190 -10 -2174
rect 52 -1798 86 -1782
rect 52 -2190 86 -2174
rect 148 -1798 182 -1782
rect 148 -2190 182 -2174
rect 244 -1798 278 -1782
rect 244 -2190 278 -2174
rect 340 -1798 374 -1782
rect 340 -2190 374 -2174
rect 436 -1798 470 -1782
rect 436 -2190 470 -2174
rect 532 -1798 566 -1782
rect 532 -2190 566 -2174
rect 628 -1798 662 -1782
rect 628 -2190 662 -2174
rect 724 -1798 758 -1782
rect 724 -2190 758 -2174
rect 820 -1798 854 -1782
rect 820 -2190 854 -2174
rect 916 -1798 950 -1782
rect 916 -2190 950 -2174
rect 1012 -1798 1046 -1782
rect 1012 -2190 1046 -2174
rect 1108 -1798 1142 -1782
rect 1108 -2190 1142 -2174
rect 1204 -1798 1238 -1782
rect 1204 -2190 1238 -2174
rect 1352 -1762 1534 -1708
rect 1352 -2070 1500 -1762
rect -1068 -2258 -1052 -2224
rect -1018 -2258 -1002 -2224
rect -876 -2258 -860 -2224
rect -826 -2258 -810 -2224
rect -684 -2258 -668 -2224
rect -634 -2258 -618 -2224
rect -492 -2258 -476 -2224
rect -442 -2258 -426 -2224
rect -300 -2258 -284 -2224
rect -250 -2258 -234 -2224
rect -108 -2258 -92 -2224
rect -58 -2258 -42 -2224
rect 84 -2258 100 -2224
rect 134 -2258 150 -2224
rect 276 -2258 292 -2224
rect 326 -2258 342 -2224
rect 468 -2258 484 -2224
rect 518 -2258 534 -2224
rect 660 -2258 676 -2224
rect 710 -2258 726 -2224
rect 852 -2258 868 -2224
rect 902 -2258 918 -2224
rect 1044 -2258 1060 -2224
rect 1094 -2258 1110 -2224
rect 1474 -2250 1500 -2070
rect -1068 -2366 -1052 -2332
rect -1018 -2366 -1002 -2332
rect -876 -2366 -860 -2332
rect -826 -2366 -810 -2332
rect -684 -2366 -668 -2332
rect -634 -2366 -618 -2332
rect -492 -2366 -476 -2332
rect -442 -2366 -426 -2332
rect -300 -2366 -284 -2332
rect -250 -2366 -234 -2332
rect -108 -2366 -92 -2332
rect -58 -2366 -42 -2332
rect 84 -2366 100 -2332
rect 134 -2366 150 -2332
rect 276 -2366 292 -2332
rect 326 -2366 342 -2332
rect 468 -2366 484 -2332
rect 518 -2366 534 -2332
rect 660 -2366 676 -2332
rect 710 -2366 726 -2332
rect 852 -2366 868 -2332
rect 902 -2366 918 -2332
rect 1044 -2366 1060 -2332
rect 1094 -2366 1110 -2332
rect -1196 -2416 -1162 -2400
rect -1196 -2808 -1162 -2792
rect -1100 -2416 -1066 -2400
rect -1100 -2808 -1066 -2792
rect -1004 -2416 -970 -2400
rect -1004 -2808 -970 -2792
rect -908 -2416 -874 -2400
rect -908 -2808 -874 -2792
rect -812 -2416 -778 -2400
rect -812 -2808 -778 -2792
rect -716 -2416 -682 -2400
rect -716 -2808 -682 -2792
rect -620 -2416 -586 -2400
rect -620 -2808 -586 -2792
rect -524 -2416 -490 -2400
rect -524 -2808 -490 -2792
rect -428 -2416 -394 -2400
rect -428 -2808 -394 -2792
rect -332 -2416 -298 -2400
rect -332 -2808 -298 -2792
rect -236 -2416 -202 -2400
rect -236 -2808 -202 -2792
rect -140 -2416 -106 -2400
rect -140 -2808 -106 -2792
rect -44 -2416 -10 -2400
rect -44 -2808 -10 -2792
rect 52 -2416 86 -2400
rect 52 -2808 86 -2792
rect 148 -2416 182 -2400
rect 148 -2808 182 -2792
rect 244 -2416 278 -2400
rect 244 -2808 278 -2792
rect 340 -2416 374 -2400
rect 340 -2808 374 -2792
rect 436 -2416 470 -2400
rect 436 -2808 470 -2792
rect 532 -2416 566 -2400
rect 532 -2808 566 -2792
rect 628 -2416 662 -2400
rect 628 -2808 662 -2792
rect 724 -2416 758 -2400
rect 724 -2808 758 -2792
rect 820 -2416 854 -2400
rect 820 -2808 854 -2792
rect 916 -2416 950 -2400
rect 916 -2808 950 -2792
rect 1012 -2416 1046 -2400
rect 1012 -2808 1046 -2792
rect 1108 -2416 1142 -2400
rect 1108 -2808 1142 -2792
rect 1204 -2416 1238 -2400
rect 1204 -2808 1238 -2792
rect -1164 -2876 -1148 -2842
rect -1114 -2876 -1098 -2842
rect -972 -2876 -956 -2842
rect -922 -2876 -906 -2842
rect -780 -2876 -764 -2842
rect -730 -2876 -714 -2842
rect -588 -2876 -572 -2842
rect -538 -2876 -522 -2842
rect -396 -2876 -380 -2842
rect -346 -2876 -330 -2842
rect -204 -2876 -188 -2842
rect -154 -2876 -138 -2842
rect -12 -2876 4 -2842
rect 38 -2876 54 -2842
rect 180 -2876 196 -2842
rect 230 -2876 246 -2842
rect 372 -2876 388 -2842
rect 422 -2876 438 -2842
rect 564 -2876 580 -2842
rect 614 -2876 630 -2842
rect 756 -2876 772 -2842
rect 806 -2876 822 -2842
rect 948 -2876 964 -2842
rect 998 -2876 1014 -2842
rect 1140 -2876 1156 -2842
rect 1190 -2876 1206 -2842
rect -1164 -2984 -1148 -2950
rect -1114 -2984 -1098 -2950
rect -972 -2984 -956 -2950
rect -922 -2984 -906 -2950
rect -780 -2984 -764 -2950
rect -730 -2984 -714 -2950
rect -588 -2984 -572 -2950
rect -538 -2984 -522 -2950
rect -396 -2984 -380 -2950
rect -346 -2984 -330 -2950
rect -204 -2984 -188 -2950
rect -154 -2984 -138 -2950
rect -12 -2984 4 -2950
rect 38 -2984 54 -2950
rect 180 -2984 196 -2950
rect 230 -2984 246 -2950
rect 372 -2984 388 -2950
rect 422 -2984 438 -2950
rect 564 -2984 580 -2950
rect 614 -2984 630 -2950
rect 756 -2984 772 -2950
rect 806 -2984 822 -2950
rect 948 -2984 964 -2950
rect 998 -2984 1014 -2950
rect 1140 -2984 1156 -2950
rect 1190 -2984 1206 -2950
rect -1196 -3034 -1162 -3018
rect -1196 -3426 -1162 -3410
rect -1100 -3034 -1066 -3018
rect -1100 -3426 -1066 -3410
rect -1004 -3034 -970 -3018
rect -1004 -3426 -970 -3410
rect -908 -3034 -874 -3018
rect -908 -3426 -874 -3410
rect -812 -3034 -778 -3018
rect -812 -3426 -778 -3410
rect -716 -3034 -682 -3018
rect -716 -3426 -682 -3410
rect -620 -3034 -586 -3018
rect -620 -3426 -586 -3410
rect -524 -3034 -490 -3018
rect -524 -3426 -490 -3410
rect -428 -3034 -394 -3018
rect -428 -3426 -394 -3410
rect -332 -3034 -298 -3018
rect -332 -3426 -298 -3410
rect -236 -3034 -202 -3018
rect -236 -3426 -202 -3410
rect -140 -3034 -106 -3018
rect -140 -3426 -106 -3410
rect -44 -3034 -10 -3018
rect -44 -3426 -10 -3410
rect 52 -3034 86 -3018
rect 52 -3426 86 -3410
rect 148 -3034 182 -3018
rect 148 -3426 182 -3410
rect 244 -3034 278 -3018
rect 244 -3426 278 -3410
rect 340 -3034 374 -3018
rect 340 -3426 374 -3410
rect 436 -3034 470 -3018
rect 436 -3426 470 -3410
rect 532 -3034 566 -3018
rect 532 -3426 566 -3410
rect 628 -3034 662 -3018
rect 628 -3426 662 -3410
rect 724 -3034 758 -3018
rect 724 -3426 758 -3410
rect 820 -3034 854 -3018
rect 820 -3426 854 -3410
rect 916 -3034 950 -3018
rect 916 -3426 950 -3410
rect 1012 -3034 1046 -3018
rect 1012 -3426 1046 -3410
rect 1108 -3034 1142 -3018
rect 1108 -3426 1142 -3410
rect 1204 -3034 1238 -3018
rect 1204 -3426 1238 -3410
rect -1068 -3494 -1052 -3460
rect -1018 -3494 -1002 -3460
rect -876 -3494 -860 -3460
rect -826 -3494 -810 -3460
rect -684 -3494 -668 -3460
rect -634 -3494 -618 -3460
rect -492 -3494 -476 -3460
rect -442 -3494 -426 -3460
rect -300 -3494 -284 -3460
rect -250 -3494 -234 -3460
rect -108 -3494 -92 -3460
rect -58 -3494 -42 -3460
rect 84 -3494 100 -3460
rect 134 -3494 150 -3460
rect 276 -3494 292 -3460
rect 326 -3494 342 -3460
rect 468 -3494 484 -3460
rect 518 -3494 534 -3460
rect 660 -3494 676 -3460
rect 710 -3494 726 -3460
rect 852 -3494 868 -3460
rect 902 -3494 918 -3460
rect 1044 -3494 1060 -3460
rect 1094 -3494 1110 -3460
rect -1068 -3602 -1052 -3568
rect -1018 -3602 -1002 -3568
rect -876 -3602 -860 -3568
rect -826 -3602 -810 -3568
rect -684 -3602 -668 -3568
rect -634 -3602 -618 -3568
rect -492 -3602 -476 -3568
rect -442 -3602 -426 -3568
rect -300 -3602 -284 -3568
rect -250 -3602 -234 -3568
rect -108 -3602 -92 -3568
rect -58 -3602 -42 -3568
rect 84 -3602 100 -3568
rect 134 -3602 150 -3568
rect 276 -3602 292 -3568
rect 326 -3602 342 -3568
rect 468 -3602 484 -3568
rect 518 -3602 534 -3568
rect 660 -3602 676 -3568
rect 710 -3602 726 -3568
rect 852 -3602 868 -3568
rect 902 -3602 918 -3568
rect 1044 -3602 1060 -3568
rect 1094 -3602 1110 -3568
rect -1196 -3652 -1162 -3636
rect -1196 -4044 -1162 -4028
rect -1100 -3652 -1066 -3636
rect -1100 -4044 -1066 -4028
rect -1004 -3652 -970 -3636
rect -1004 -4044 -970 -4028
rect -908 -3652 -874 -3636
rect -908 -4044 -874 -4028
rect -812 -3652 -778 -3636
rect -812 -4044 -778 -4028
rect -716 -3652 -682 -3636
rect -716 -4044 -682 -4028
rect -620 -3652 -586 -3636
rect -620 -4044 -586 -4028
rect -524 -3652 -490 -3636
rect -524 -4044 -490 -4028
rect -428 -3652 -394 -3636
rect -428 -4044 -394 -4028
rect -332 -3652 -298 -3636
rect -332 -4044 -298 -4028
rect -236 -3652 -202 -3636
rect -236 -4044 -202 -4028
rect -140 -3652 -106 -3636
rect -140 -4044 -106 -4028
rect -44 -3652 -10 -3636
rect -44 -4044 -10 -4028
rect 52 -3652 86 -3636
rect 52 -4044 86 -4028
rect 148 -3652 182 -3636
rect 148 -4044 182 -4028
rect 244 -3652 278 -3636
rect 244 -4044 278 -4028
rect 340 -3652 374 -3636
rect 340 -4044 374 -4028
rect 436 -3652 470 -3636
rect 436 -4044 470 -4028
rect 532 -3652 566 -3636
rect 532 -4044 566 -4028
rect 628 -3652 662 -3636
rect 628 -4044 662 -4028
rect 724 -3652 758 -3636
rect 724 -4044 758 -4028
rect 820 -3652 854 -3636
rect 820 -4044 854 -4028
rect 916 -3652 950 -3636
rect 916 -4044 950 -4028
rect 1012 -3652 1046 -3636
rect 1012 -4044 1046 -4028
rect 1108 -3652 1142 -3636
rect 1108 -4044 1142 -4028
rect 1204 -3652 1238 -3636
rect 1204 -4044 1238 -4028
rect -1164 -4112 -1148 -4078
rect -1114 -4112 -1098 -4078
rect -972 -4112 -956 -4078
rect -922 -4112 -906 -4078
rect -780 -4112 -764 -4078
rect -730 -4112 -714 -4078
rect -588 -4112 -572 -4078
rect -538 -4112 -522 -4078
rect -396 -4112 -380 -4078
rect -346 -4112 -330 -4078
rect -204 -4112 -188 -4078
rect -154 -4112 -138 -4078
rect -12 -4112 4 -4078
rect 38 -4112 54 -4078
rect 180 -4112 196 -4078
rect 230 -4112 246 -4078
rect 372 -4112 388 -4078
rect 422 -4112 438 -4078
rect 564 -4112 580 -4078
rect 614 -4112 630 -4078
rect 756 -4112 772 -4078
rect 806 -4112 822 -4078
rect 948 -4112 964 -4078
rect 998 -4112 1014 -4078
rect 1140 -4112 1156 -4078
rect 1190 -4112 1206 -4078
rect -1396 -4180 -1256 -4118
rect 1352 -2318 1500 -2250
rect 3276 -1762 3310 -1700
rect 1660 -1802 1676 -1768
rect 1844 -1802 1860 -1768
rect 1918 -1802 1934 -1768
rect 2102 -1802 2118 -1768
rect 2176 -1802 2192 -1768
rect 2360 -1802 2376 -1768
rect 2434 -1802 2450 -1768
rect 2618 -1802 2634 -1768
rect 2692 -1802 2708 -1768
rect 2876 -1802 2892 -1768
rect 2950 -1802 2966 -1768
rect 3134 -1802 3150 -1768
rect 1614 -1852 1648 -1836
rect 1614 -2244 1648 -2228
rect 1872 -1852 1906 -1836
rect 1872 -2244 1906 -2228
rect 2130 -1852 2164 -1836
rect 2130 -2244 2164 -2228
rect 2388 -1852 2422 -1836
rect 2388 -2244 2422 -2228
rect 2646 -1852 2680 -1836
rect 2646 -2244 2680 -2228
rect 2904 -1852 2938 -1836
rect 2904 -2244 2938 -2228
rect 3162 -1852 3196 -1836
rect 3162 -2244 3196 -2228
rect 1660 -2312 1676 -2278
rect 1844 -2312 1860 -2278
rect 1918 -2312 1934 -2278
rect 2102 -2312 2118 -2278
rect 2176 -2312 2192 -2278
rect 2360 -2312 2376 -2278
rect 2434 -2312 2450 -2278
rect 2618 -2312 2634 -2278
rect 2692 -2312 2708 -2278
rect 2876 -2312 2892 -2278
rect 2950 -2312 2966 -2278
rect 3134 -2312 3150 -2278
rect 1352 -2380 1534 -2318
rect 3230 -2318 3276 -2130
rect 3310 -2318 5340 -2130
rect 3230 -2380 5340 -2318
rect 1352 -2414 1596 -2380
rect 3214 -2414 5340 -2380
rect 1352 -2570 5340 -2414
rect 1318 -4180 1352 -4118
rect -1396 -4214 -1214 -4180
rect 1256 -4214 1352 -4180
rect -1396 -4220 -1256 -4214
rect -1296 -4342 2324 -4280
rect -1296 -4360 -1194 -4342
rect -1290 -4376 -1194 -4360
rect 346 -4376 604 -4342
rect 2144 -4376 2324 -4342
rect -1290 -4438 -1256 -4376
rect 408 -4438 542 -4376
rect -1143 -4478 -1127 -4444
rect -1093 -4478 -1029 -4444
rect -995 -4478 -931 -4444
rect -897 -4478 -833 -4444
rect -799 -4478 -735 -4444
rect -701 -4478 -637 -4444
rect -603 -4478 -539 -4444
rect -505 -4478 -441 -4444
rect -407 -4478 -343 -4444
rect -309 -4478 -245 -4444
rect -211 -4478 -147 -4444
rect -113 -4478 -49 -4444
rect -15 -4478 49 -4444
rect 83 -4478 147 -4444
rect 181 -4478 245 -4444
rect 279 -4478 295 -4444
rect -1176 -4537 -1142 -4521
rect -1176 -4929 -1142 -4913
rect -1078 -4537 -1044 -4521
rect -1078 -4929 -1044 -4913
rect -980 -4537 -946 -4521
rect -980 -4929 -946 -4913
rect -882 -4537 -848 -4521
rect -882 -4929 -848 -4913
rect -784 -4537 -750 -4521
rect -784 -4929 -750 -4913
rect -686 -4537 -652 -4521
rect -686 -4929 -652 -4913
rect -588 -4537 -554 -4521
rect -588 -4929 -554 -4913
rect -490 -4537 -456 -4521
rect -490 -4929 -456 -4913
rect -392 -4537 -358 -4521
rect -392 -4929 -358 -4913
rect -294 -4537 -260 -4521
rect -294 -4929 -260 -4913
rect -196 -4537 -162 -4521
rect -196 -4929 -162 -4913
rect -98 -4537 -64 -4521
rect -98 -4929 -64 -4913
rect 0 -4537 34 -4521
rect 0 -4929 34 -4913
rect 98 -4537 132 -4521
rect 98 -4929 132 -4913
rect 196 -4537 230 -4521
rect 196 -4929 230 -4913
rect 294 -4537 328 -4521
rect 294 -4929 328 -4913
rect -1143 -5006 -1127 -4972
rect -1093 -5006 -1029 -4972
rect -995 -5006 -931 -4972
rect -897 -5006 -833 -4972
rect -799 -5006 -735 -4972
rect -701 -5006 -637 -4972
rect -603 -5006 -539 -4972
rect -505 -5006 -441 -4972
rect -407 -5006 -343 -4972
rect -309 -5006 -245 -4972
rect -211 -5006 -147 -4972
rect -113 -5006 -49 -4972
rect -15 -5006 49 -4972
rect 83 -5006 147 -4972
rect 181 -5006 245 -4972
rect 279 -5006 295 -4972
rect -1143 -5114 -1127 -5080
rect -1093 -5114 -1029 -5080
rect -995 -5114 -931 -5080
rect -897 -5114 -833 -5080
rect -799 -5114 -735 -5080
rect -701 -5114 -637 -5080
rect -603 -5114 -539 -5080
rect -505 -5114 -441 -5080
rect -407 -5114 -343 -5080
rect -309 -5114 -245 -5080
rect -211 -5114 -147 -5080
rect -113 -5114 -49 -5080
rect -15 -5114 49 -5080
rect 83 -5114 147 -5080
rect 181 -5114 245 -5080
rect 279 -5114 295 -5080
rect -1176 -5173 -1142 -5157
rect -1176 -5565 -1142 -5549
rect -1078 -5173 -1044 -5157
rect -1078 -5565 -1044 -5549
rect -980 -5173 -946 -5157
rect -980 -5565 -946 -5549
rect -882 -5173 -848 -5157
rect -882 -5565 -848 -5549
rect -784 -5173 -750 -5157
rect -784 -5565 -750 -5549
rect -686 -5173 -652 -5157
rect -686 -5565 -652 -5549
rect -588 -5173 -554 -5157
rect -588 -5565 -554 -5549
rect -490 -5173 -456 -5157
rect -490 -5565 -456 -5549
rect -392 -5173 -358 -5157
rect -392 -5565 -358 -5549
rect -294 -5173 -260 -5157
rect -294 -5565 -260 -5549
rect -196 -5173 -162 -5157
rect -196 -5565 -162 -5549
rect -98 -5173 -64 -5157
rect -98 -5565 -64 -5549
rect 0 -5173 34 -5157
rect 0 -5565 34 -5549
rect 98 -5173 132 -5157
rect 98 -5565 132 -5549
rect 196 -5173 230 -5157
rect 196 -5565 230 -5549
rect 294 -5173 328 -5157
rect 294 -5565 328 -5549
rect -1143 -5642 -1127 -5608
rect -1093 -5642 -1029 -5608
rect -995 -5642 -931 -5608
rect -897 -5642 -833 -5608
rect -799 -5642 -735 -5608
rect -701 -5642 -637 -5608
rect -603 -5642 -539 -5608
rect -505 -5642 -441 -5608
rect -407 -5642 -343 -5608
rect -309 -5642 -245 -5608
rect -211 -5642 -147 -5608
rect -113 -5642 -49 -5608
rect -15 -5642 49 -5608
rect 83 -5642 147 -5608
rect 181 -5642 245 -5608
rect 279 -5642 295 -5608
rect -1290 -5710 -1256 -5648
rect 442 -5648 508 -4438
rect 2206 -4438 2324 -4376
rect 655 -4478 671 -4444
rect 705 -4478 769 -4444
rect 803 -4478 867 -4444
rect 901 -4478 965 -4444
rect 999 -4478 1063 -4444
rect 1097 -4478 1161 -4444
rect 1195 -4478 1259 -4444
rect 1293 -4478 1357 -4444
rect 1391 -4478 1455 -4444
rect 1489 -4478 1553 -4444
rect 1587 -4478 1651 -4444
rect 1685 -4478 1749 -4444
rect 1783 -4478 1847 -4444
rect 1881 -4478 1945 -4444
rect 1979 -4478 2043 -4444
rect 2077 -4478 2093 -4444
rect 622 -4537 656 -4521
rect 622 -4929 656 -4913
rect 720 -4537 754 -4521
rect 720 -4929 754 -4913
rect 818 -4537 852 -4521
rect 818 -4929 852 -4913
rect 916 -4537 950 -4521
rect 916 -4929 950 -4913
rect 1014 -4537 1048 -4521
rect 1014 -4929 1048 -4913
rect 1112 -4537 1146 -4521
rect 1112 -4929 1146 -4913
rect 1210 -4537 1244 -4521
rect 1210 -4929 1244 -4913
rect 1308 -4537 1342 -4521
rect 1308 -4929 1342 -4913
rect 1406 -4537 1440 -4521
rect 1406 -4929 1440 -4913
rect 1504 -4537 1538 -4521
rect 1504 -4929 1538 -4913
rect 1602 -4537 1636 -4521
rect 1602 -4929 1636 -4913
rect 1700 -4537 1734 -4521
rect 1700 -4929 1734 -4913
rect 1798 -4537 1832 -4521
rect 1798 -4929 1832 -4913
rect 1896 -4537 1930 -4521
rect 1896 -4929 1930 -4913
rect 1994 -4537 2028 -4521
rect 1994 -4929 2028 -4913
rect 2092 -4537 2126 -4521
rect 2092 -4929 2126 -4913
rect 655 -5006 671 -4972
rect 705 -5006 769 -4972
rect 803 -5006 867 -4972
rect 901 -5006 965 -4972
rect 999 -5006 1063 -4972
rect 1097 -5006 1161 -4972
rect 1195 -5006 1259 -4972
rect 1293 -5006 1357 -4972
rect 1391 -5006 1455 -4972
rect 1489 -5006 1553 -4972
rect 1587 -5006 1651 -4972
rect 1685 -5006 1749 -4972
rect 1783 -5006 1847 -4972
rect 1881 -5006 1945 -4972
rect 1979 -5006 2043 -4972
rect 2077 -5006 2093 -4972
rect 2240 -4910 2324 -4438
rect 2240 -4994 4394 -4910
rect 2240 -5000 2406 -4994
rect 655 -5114 671 -5080
rect 705 -5114 769 -5080
rect 803 -5114 867 -5080
rect 901 -5114 965 -5080
rect 999 -5114 1063 -5080
rect 1097 -5114 1161 -5080
rect 1195 -5114 1259 -5080
rect 1293 -5114 1357 -5080
rect 1391 -5114 1455 -5080
rect 1489 -5114 1553 -5080
rect 1587 -5114 1651 -5080
rect 1685 -5114 1749 -5080
rect 1783 -5114 1847 -5080
rect 1881 -5114 1945 -5080
rect 1979 -5114 2043 -5080
rect 2077 -5114 2093 -5080
rect 622 -5173 656 -5157
rect 622 -5565 656 -5549
rect 720 -5173 754 -5157
rect 720 -5565 754 -5549
rect 818 -5173 852 -5157
rect 818 -5565 852 -5549
rect 916 -5173 950 -5157
rect 916 -5565 950 -5549
rect 1014 -5173 1048 -5157
rect 1014 -5565 1048 -5549
rect 1112 -5173 1146 -5157
rect 1112 -5565 1146 -5549
rect 1210 -5173 1244 -5157
rect 1210 -5565 1244 -5549
rect 1308 -5173 1342 -5157
rect 1308 -5565 1342 -5549
rect 1406 -5173 1440 -5157
rect 1406 -5565 1440 -5549
rect 1504 -5173 1538 -5157
rect 1504 -5565 1538 -5549
rect 1602 -5173 1636 -5157
rect 1602 -5565 1636 -5549
rect 1700 -5173 1734 -5157
rect 1700 -5565 1734 -5549
rect 1798 -5173 1832 -5157
rect 1798 -5565 1832 -5549
rect 1896 -5173 1930 -5157
rect 1896 -5565 1930 -5549
rect 1994 -5173 2028 -5157
rect 1994 -5565 2028 -5549
rect 2092 -5173 2126 -5157
rect 2092 -5565 2126 -5549
rect 2344 -5028 2406 -5000
rect 4056 -5028 4394 -4994
rect 4118 -5090 4394 -5028
rect 2470 -5130 2486 -5096
rect 2554 -5130 2570 -5096
rect 2628 -5130 2644 -5096
rect 2712 -5130 2728 -5096
rect 2786 -5130 2802 -5096
rect 2870 -5130 2886 -5096
rect 2944 -5130 2960 -5096
rect 3028 -5130 3044 -5096
rect 3102 -5130 3118 -5096
rect 3186 -5130 3202 -5096
rect 3260 -5130 3276 -5096
rect 3344 -5130 3360 -5096
rect 3418 -5130 3434 -5096
rect 3502 -5130 3518 -5096
rect 3576 -5130 3592 -5096
rect 3660 -5130 3676 -5096
rect 3734 -5130 3750 -5096
rect 3818 -5130 3834 -5096
rect 3892 -5130 3908 -5096
rect 3976 -5130 3992 -5096
rect 655 -5642 671 -5608
rect 705 -5642 769 -5608
rect 803 -5642 867 -5608
rect 901 -5642 965 -5608
rect 999 -5642 1063 -5608
rect 1097 -5642 1161 -5608
rect 1195 -5642 1259 -5608
rect 1293 -5642 1357 -5608
rect 1391 -5642 1455 -5608
rect 1489 -5642 1553 -5608
rect 1587 -5642 1651 -5608
rect 1685 -5642 1749 -5608
rect 1783 -5642 1847 -5608
rect 1881 -5642 1945 -5608
rect 1979 -5642 2043 -5608
rect 2077 -5642 2093 -5608
rect 408 -5710 542 -5648
rect 2240 -5648 2310 -5560
rect 2206 -5664 2310 -5648
rect 2424 -5189 2458 -5173
rect 2424 -5581 2458 -5565
rect 2582 -5189 2616 -5173
rect 2582 -5581 2616 -5565
rect 2740 -5189 2774 -5173
rect 2740 -5581 2774 -5565
rect 2898 -5189 2932 -5173
rect 2898 -5581 2932 -5565
rect 3056 -5189 3090 -5173
rect 3056 -5581 3090 -5565
rect 3214 -5189 3248 -5173
rect 3214 -5581 3248 -5565
rect 3372 -5189 3406 -5173
rect 3372 -5581 3406 -5565
rect 3530 -5189 3564 -5173
rect 3530 -5581 3564 -5565
rect 3688 -5189 3722 -5173
rect 3688 -5581 3722 -5565
rect 3846 -5189 3880 -5173
rect 3846 -5581 3880 -5565
rect 4004 -5189 4038 -5173
rect 4004 -5581 4038 -5565
rect 2470 -5658 2486 -5624
rect 2554 -5658 2570 -5624
rect 2628 -5658 2644 -5624
rect 2712 -5658 2728 -5624
rect 2786 -5658 2802 -5624
rect 2870 -5658 2886 -5624
rect 2944 -5658 2960 -5624
rect 3028 -5658 3044 -5624
rect 3102 -5658 3118 -5624
rect 3186 -5658 3202 -5624
rect 3260 -5658 3276 -5624
rect 3344 -5658 3360 -5624
rect 3418 -5658 3434 -5624
rect 3502 -5658 3518 -5624
rect 3576 -5658 3592 -5624
rect 3660 -5658 3676 -5624
rect 3734 -5658 3750 -5624
rect 3818 -5658 3834 -5624
rect 3892 -5658 3908 -5624
rect 3976 -5658 3992 -5624
rect 2206 -5710 2344 -5664
rect -1290 -5744 -1194 -5710
rect 346 -5740 604 -5710
rect 346 -5744 442 -5740
rect 508 -5744 604 -5740
rect 2144 -5726 2344 -5710
rect 4152 -5664 4394 -5090
rect 4118 -5726 4394 -5664
rect 2144 -5744 2406 -5726
rect 2074 -5760 2406 -5744
rect 4056 -5760 4394 -5726
rect -1290 -5830 -1194 -5818
rect -1396 -5852 -1194 -5830
rect 1326 -5820 1422 -5818
rect 1326 -5852 1534 -5820
rect 2074 -5837 4394 -5760
rect -1396 -5914 -1256 -5852
rect -1396 -7088 -1290 -5914
rect 1388 -5914 1534 -5852
rect -1144 -5954 -1127 -5920
rect -1093 -5954 -1030 -5920
rect -996 -5954 -931 -5920
rect -897 -5954 -834 -5920
rect -800 -5954 -735 -5920
rect -701 -5954 -638 -5920
rect -604 -5954 -539 -5920
rect -505 -5954 -442 -5920
rect -408 -5954 -343 -5920
rect -309 -5954 -246 -5920
rect -212 -5954 -147 -5920
rect -113 -5954 -50 -5920
rect -16 -5954 49 -5920
rect 83 -5954 146 -5920
rect 180 -5954 245 -5920
rect 279 -5954 342 -5920
rect 376 -5954 441 -5920
rect 475 -5954 538 -5920
rect 572 -5954 637 -5920
rect 671 -5954 734 -5920
rect 768 -5954 833 -5920
rect 867 -5954 930 -5920
rect 964 -5954 1029 -5920
rect 1063 -5954 1126 -5920
rect 1160 -5954 1225 -5920
rect 1259 -5954 1275 -5920
rect -1176 -6004 -1142 -5988
rect -1176 -6396 -1142 -6380
rect -1078 -6004 -1044 -5988
rect -1078 -6396 -1044 -6380
rect -980 -6004 -946 -5988
rect -980 -6396 -946 -6380
rect -882 -6004 -848 -5988
rect -882 -6396 -848 -6380
rect -784 -6004 -750 -5988
rect -784 -6396 -750 -6380
rect -686 -6004 -652 -5988
rect -686 -6396 -652 -6380
rect -588 -6004 -554 -5988
rect -588 -6396 -554 -6380
rect -490 -6004 -456 -5988
rect -490 -6396 -456 -6380
rect -392 -6004 -358 -5988
rect -392 -6396 -358 -6380
rect -294 -6004 -260 -5988
rect -294 -6396 -260 -6380
rect -196 -6004 -162 -5988
rect -196 -6396 -162 -6380
rect -98 -6004 -64 -5988
rect -98 -6396 -64 -6380
rect 0 -6004 34 -5988
rect 0 -6396 34 -6380
rect 98 -6004 132 -5988
rect 98 -6396 132 -6380
rect 196 -6004 230 -5988
rect 196 -6396 230 -6380
rect 294 -6004 328 -5988
rect 294 -6396 328 -6380
rect 392 -6004 426 -5988
rect 392 -6396 426 -6380
rect 490 -6004 524 -5988
rect 490 -6396 524 -6380
rect 588 -6004 622 -5988
rect 588 -6396 622 -6380
rect 686 -6004 720 -5988
rect 686 -6396 720 -6380
rect 784 -6004 818 -5988
rect 784 -6396 818 -6380
rect 882 -6004 916 -5988
rect 882 -6396 916 -6380
rect 980 -6004 1014 -5988
rect 980 -6396 1014 -6380
rect 1078 -6004 1112 -5988
rect 1078 -6396 1112 -6380
rect 1176 -6004 1210 -5988
rect 1176 -6396 1210 -6380
rect 1274 -6004 1308 -5988
rect 1274 -6396 1308 -6380
rect -1144 -6464 -1128 -6430
rect -1094 -6464 -1029 -6430
rect -995 -6464 -932 -6430
rect -898 -6464 -833 -6430
rect -799 -6464 -736 -6430
rect -702 -6464 -637 -6430
rect -603 -6464 -540 -6430
rect -506 -6464 -441 -6430
rect -407 -6464 -344 -6430
rect -310 -6464 -245 -6430
rect -211 -6464 -148 -6430
rect -114 -6464 -49 -6430
rect -15 -6464 48 -6430
rect 82 -6464 147 -6430
rect 181 -6464 244 -6430
rect 278 -6464 343 -6430
rect 377 -6464 440 -6430
rect 474 -6464 539 -6430
rect 573 -6464 636 -6430
rect 670 -6464 735 -6430
rect 769 -6464 832 -6430
rect 866 -6464 931 -6430
rect 965 -6464 1028 -6430
rect 1062 -6464 1127 -6430
rect 1161 -6464 1224 -6430
rect 1258 -6464 1274 -6430
rect -1143 -6572 -1127 -6538
rect -1093 -6572 -1029 -6538
rect -995 -6572 -931 -6538
rect -897 -6572 -833 -6538
rect -799 -6572 -735 -6538
rect -701 -6572 -637 -6538
rect -603 -6572 -539 -6538
rect -505 -6572 -441 -6538
rect -407 -6572 -343 -6538
rect -309 -6572 -245 -6538
rect -211 -6572 -147 -6538
rect -113 -6572 -49 -6538
rect -15 -6572 49 -6538
rect 83 -6572 147 -6538
rect 181 -6572 245 -6538
rect 279 -6572 343 -6538
rect 377 -6572 441 -6538
rect 475 -6572 539 -6538
rect 573 -6572 637 -6538
rect 671 -6572 735 -6538
rect 769 -6572 833 -6538
rect 867 -6572 931 -6538
rect 965 -6572 1029 -6538
rect 1063 -6572 1127 -6538
rect 1161 -6572 1225 -6538
rect 1259 -6572 1275 -6538
rect -1176 -6622 -1142 -6606
rect -1176 -7014 -1142 -6998
rect -1078 -6622 -1044 -6606
rect -1078 -7014 -1044 -6998
rect -980 -6622 -946 -6606
rect -980 -7014 -946 -6998
rect -882 -6622 -848 -6606
rect -882 -7014 -848 -6998
rect -784 -6622 -750 -6606
rect -784 -7014 -750 -6998
rect -686 -6622 -652 -6606
rect -686 -7014 -652 -6998
rect -588 -6622 -554 -6606
rect -588 -7014 -554 -6998
rect -490 -6622 -456 -6606
rect -490 -7014 -456 -6998
rect -392 -6622 -358 -6606
rect -392 -7014 -358 -6998
rect -294 -6622 -260 -6606
rect -294 -7014 -260 -6998
rect -196 -6622 -162 -6606
rect -196 -7014 -162 -6998
rect -98 -6622 -64 -6606
rect -98 -7014 -64 -6998
rect 0 -6622 34 -6606
rect 0 -7014 34 -6998
rect 98 -6622 132 -6606
rect 98 -7014 132 -6998
rect 196 -6622 230 -6606
rect 196 -7014 230 -6998
rect 294 -6622 328 -6606
rect 294 -7014 328 -6998
rect 392 -6622 426 -6606
rect 392 -7014 426 -6998
rect 490 -6622 524 -6606
rect 490 -7014 524 -6998
rect 588 -6622 622 -6606
rect 588 -7014 622 -6998
rect 686 -6622 720 -6606
rect 686 -7014 720 -6998
rect 784 -6622 818 -6606
rect 784 -7014 818 -6998
rect 882 -6622 916 -6606
rect 882 -7014 916 -6998
rect 980 -6622 1014 -6606
rect 980 -7014 1014 -6998
rect 1078 -6622 1112 -6606
rect 1078 -7014 1112 -6998
rect 1176 -6622 1210 -6606
rect 1176 -7014 1210 -6998
rect 1274 -6622 1308 -6606
rect 1274 -7014 1308 -6998
rect -1143 -7082 -1127 -7048
rect -1093 -7082 -1029 -7048
rect -995 -7082 -931 -7048
rect -897 -7082 -833 -7048
rect -799 -7082 -735 -7048
rect -701 -7082 -637 -7048
rect -603 -7082 -539 -7048
rect -505 -7082 -441 -7048
rect -407 -7082 -343 -7048
rect -309 -7082 -245 -7048
rect -211 -7082 -147 -7048
rect -113 -7082 -49 -7048
rect -15 -7082 49 -7048
rect 83 -7082 147 -7048
rect 181 -7082 245 -7048
rect 279 -7082 343 -7048
rect 377 -7082 441 -7048
rect 475 -7082 539 -7048
rect 573 -7082 637 -7048
rect 671 -7082 735 -7048
rect 769 -7082 833 -7048
rect 867 -7082 931 -7048
rect 965 -7082 1029 -7048
rect 1063 -7082 1127 -7048
rect 1161 -7082 1225 -7048
rect 1259 -7082 1275 -7048
rect -1396 -7150 -1256 -7088
rect 1422 -7088 1534 -5914
rect 1388 -7150 1534 -7088
rect -1396 -7184 -1194 -7150
rect 1326 -7184 1534 -7150
rect -1396 -7262 1534 -7184
rect -1396 -7296 -1194 -7262
rect 1326 -7296 1534 -7262
rect -1396 -7358 -1256 -7296
rect -1396 -8532 -1290 -7358
rect 1388 -7358 1534 -7296
rect -1144 -7398 -1127 -7364
rect -1093 -7398 -1030 -7364
rect -996 -7398 -931 -7364
rect -897 -7398 -834 -7364
rect -800 -7398 -735 -7364
rect -701 -7398 -638 -7364
rect -604 -7398 -539 -7364
rect -505 -7398 -442 -7364
rect -408 -7398 -343 -7364
rect -309 -7398 -246 -7364
rect -212 -7398 -147 -7364
rect -113 -7398 -50 -7364
rect -16 -7398 49 -7364
rect 83 -7398 146 -7364
rect 180 -7398 245 -7364
rect 279 -7398 342 -7364
rect 376 -7398 441 -7364
rect 475 -7398 538 -7364
rect 572 -7398 637 -7364
rect 671 -7398 734 -7364
rect 768 -7398 833 -7364
rect 867 -7398 930 -7364
rect 964 -7398 1029 -7364
rect 1063 -7398 1126 -7364
rect 1160 -7398 1225 -7364
rect 1259 -7398 1275 -7364
rect -1176 -7448 -1142 -7432
rect -1176 -7840 -1142 -7824
rect -1078 -7448 -1044 -7432
rect -1078 -7840 -1044 -7824
rect -980 -7448 -946 -7432
rect -980 -7840 -946 -7824
rect -882 -7448 -848 -7432
rect -882 -7840 -848 -7824
rect -784 -7448 -750 -7432
rect -784 -7840 -750 -7824
rect -686 -7448 -652 -7432
rect -686 -7840 -652 -7824
rect -588 -7448 -554 -7432
rect -588 -7840 -554 -7824
rect -490 -7448 -456 -7432
rect -490 -7840 -456 -7824
rect -392 -7448 -358 -7432
rect -392 -7840 -358 -7824
rect -294 -7448 -260 -7432
rect -294 -7840 -260 -7824
rect -196 -7448 -162 -7432
rect -196 -7840 -162 -7824
rect -98 -7448 -64 -7432
rect -98 -7840 -64 -7824
rect 0 -7448 34 -7432
rect 0 -7840 34 -7824
rect 98 -7448 132 -7432
rect 98 -7840 132 -7824
rect 196 -7448 230 -7432
rect 196 -7840 230 -7824
rect 294 -7448 328 -7432
rect 294 -7840 328 -7824
rect 392 -7448 426 -7432
rect 392 -7840 426 -7824
rect 490 -7448 524 -7432
rect 490 -7840 524 -7824
rect 588 -7448 622 -7432
rect 588 -7840 622 -7824
rect 686 -7448 720 -7432
rect 686 -7840 720 -7824
rect 784 -7448 818 -7432
rect 784 -7840 818 -7824
rect 882 -7448 916 -7432
rect 882 -7840 916 -7824
rect 980 -7448 1014 -7432
rect 980 -7840 1014 -7824
rect 1078 -7448 1112 -7432
rect 1078 -7840 1112 -7824
rect 1176 -7448 1210 -7432
rect 1176 -7840 1210 -7824
rect 1274 -7448 1308 -7432
rect 1274 -7840 1308 -7824
rect -1144 -7908 -1128 -7874
rect -1094 -7908 -1029 -7874
rect -995 -7908 -932 -7874
rect -898 -7908 -833 -7874
rect -799 -7908 -736 -7874
rect -702 -7908 -637 -7874
rect -603 -7908 -540 -7874
rect -506 -7908 -441 -7874
rect -407 -7908 -344 -7874
rect -310 -7908 -245 -7874
rect -211 -7908 -148 -7874
rect -114 -7908 -49 -7874
rect -15 -7908 48 -7874
rect 82 -7908 147 -7874
rect 181 -7908 244 -7874
rect 278 -7908 343 -7874
rect 377 -7908 440 -7874
rect 474 -7908 539 -7874
rect 573 -7908 636 -7874
rect 670 -7908 735 -7874
rect 769 -7908 832 -7874
rect 866 -7908 931 -7874
rect 965 -7908 1028 -7874
rect 1062 -7908 1127 -7874
rect 1161 -7908 1224 -7874
rect 1258 -7908 1274 -7874
rect -1143 -8016 -1127 -7982
rect -1093 -8016 -1029 -7982
rect -995 -8016 -931 -7982
rect -897 -8016 -833 -7982
rect -799 -8016 -735 -7982
rect -701 -8016 -637 -7982
rect -603 -8016 -539 -7982
rect -505 -8016 -441 -7982
rect -407 -8016 -343 -7982
rect -309 -8016 -245 -7982
rect -211 -8016 -147 -7982
rect -113 -8016 -49 -7982
rect -15 -8016 49 -7982
rect 83 -8016 147 -7982
rect 181 -8016 245 -7982
rect 279 -8016 343 -7982
rect 377 -8016 441 -7982
rect 475 -8016 539 -7982
rect 573 -8016 637 -7982
rect 671 -8016 735 -7982
rect 769 -8016 833 -7982
rect 867 -8016 931 -7982
rect 965 -8016 1029 -7982
rect 1063 -8016 1127 -7982
rect 1161 -8016 1225 -7982
rect 1259 -8016 1275 -7982
rect -1176 -8066 -1142 -8050
rect -1176 -8458 -1142 -8442
rect -1078 -8066 -1044 -8050
rect -1078 -8458 -1044 -8442
rect -980 -8066 -946 -8050
rect -980 -8458 -946 -8442
rect -882 -8066 -848 -8050
rect -882 -8458 -848 -8442
rect -784 -8066 -750 -8050
rect -784 -8458 -750 -8442
rect -686 -8066 -652 -8050
rect -686 -8458 -652 -8442
rect -588 -8066 -554 -8050
rect -588 -8458 -554 -8442
rect -490 -8066 -456 -8050
rect -490 -8458 -456 -8442
rect -392 -8066 -358 -8050
rect -392 -8458 -358 -8442
rect -294 -8066 -260 -8050
rect -294 -8458 -260 -8442
rect -196 -8066 -162 -8050
rect -196 -8458 -162 -8442
rect -98 -8066 -64 -8050
rect -98 -8458 -64 -8442
rect 0 -8066 34 -8050
rect 0 -8458 34 -8442
rect 98 -8066 132 -8050
rect 98 -8458 132 -8442
rect 196 -8066 230 -8050
rect 196 -8458 230 -8442
rect 294 -8066 328 -8050
rect 294 -8458 328 -8442
rect 392 -8066 426 -8050
rect 392 -8458 426 -8442
rect 490 -8066 524 -8050
rect 490 -8458 524 -8442
rect 588 -8066 622 -8050
rect 588 -8458 622 -8442
rect 686 -8066 720 -8050
rect 686 -8458 720 -8442
rect 784 -8066 818 -8050
rect 784 -8458 818 -8442
rect 882 -8066 916 -8050
rect 882 -8458 916 -8442
rect 980 -8066 1014 -8050
rect 980 -8458 1014 -8442
rect 1078 -8066 1112 -8050
rect 1078 -8458 1112 -8442
rect 1176 -8066 1210 -8050
rect 1176 -8458 1210 -8442
rect 1274 -8066 1308 -8050
rect 1274 -8458 1308 -8442
rect -1143 -8526 -1127 -8492
rect -1093 -8526 -1029 -8492
rect -995 -8526 -931 -8492
rect -897 -8526 -833 -8492
rect -799 -8526 -735 -8492
rect -701 -8526 -637 -8492
rect -603 -8526 -539 -8492
rect -505 -8526 -441 -8492
rect -407 -8526 -343 -8492
rect -309 -8526 -245 -8492
rect -211 -8526 -147 -8492
rect -113 -8526 -49 -8492
rect -15 -8526 49 -8492
rect 83 -8526 147 -8492
rect 181 -8526 245 -8492
rect 279 -8526 343 -8492
rect 377 -8526 441 -8492
rect 475 -8526 539 -8492
rect 573 -8526 637 -8492
rect 671 -8526 735 -8492
rect 769 -8526 833 -8492
rect 867 -8526 931 -8492
rect 965 -8526 1029 -8492
rect 1063 -8526 1127 -8492
rect 1161 -8526 1225 -8492
rect 1259 -8526 1275 -8492
rect -1396 -8594 -1256 -8532
rect 1422 -7916 1534 -7358
rect 2071 -5871 2131 -5837
rect 4337 -5871 4397 -5837
rect 2071 -5897 2105 -5871
rect 4363 -5897 4397 -5871
rect 2304 -6138 4174 -6070
rect 2304 -6172 2466 -6138
rect 4006 -6172 4174 -6138
rect 2304 -6234 2404 -6172
rect 2304 -6750 2370 -6234
rect 2284 -6910 2370 -6750
rect 2294 -7408 2370 -6910
rect 4068 -6234 4174 -6172
rect 2517 -6274 2533 -6240
rect 2567 -6274 2631 -6240
rect 2665 -6274 2729 -6240
rect 2763 -6274 2827 -6240
rect 2861 -6274 2925 -6240
rect 2959 -6274 3023 -6240
rect 3057 -6274 3121 -6240
rect 3155 -6274 3219 -6240
rect 3253 -6274 3317 -6240
rect 3351 -6274 3415 -6240
rect 3449 -6274 3513 -6240
rect 3547 -6274 3611 -6240
rect 3645 -6274 3709 -6240
rect 3743 -6274 3807 -6240
rect 3841 -6274 3905 -6240
rect 3939 -6274 3955 -6240
rect 2484 -6324 2518 -6308
rect 2484 -6716 2518 -6700
rect 2582 -6324 2616 -6308
rect 2582 -6716 2616 -6700
rect 2680 -6324 2714 -6308
rect 2680 -6716 2714 -6700
rect 2778 -6324 2812 -6308
rect 2778 -6716 2812 -6700
rect 2876 -6324 2910 -6308
rect 2876 -6716 2910 -6700
rect 2974 -6324 3008 -6308
rect 2974 -6716 3008 -6700
rect 3072 -6324 3106 -6308
rect 3072 -6716 3106 -6700
rect 3170 -6324 3204 -6308
rect 3170 -6716 3204 -6700
rect 3268 -6324 3302 -6308
rect 3268 -6716 3302 -6700
rect 3366 -6324 3400 -6308
rect 3366 -6716 3400 -6700
rect 3464 -6324 3498 -6308
rect 3464 -6716 3498 -6700
rect 3562 -6324 3596 -6308
rect 3562 -6716 3596 -6700
rect 3660 -6324 3694 -6308
rect 3660 -6716 3694 -6700
rect 3758 -6324 3792 -6308
rect 3758 -6716 3792 -6700
rect 3856 -6324 3890 -6308
rect 3856 -6716 3890 -6700
rect 3954 -6324 3988 -6308
rect 3954 -6716 3988 -6700
rect 4102 -6730 4174 -6234
rect 2517 -6784 2533 -6750
rect 2567 -6784 2631 -6750
rect 2665 -6784 2729 -6750
rect 2763 -6784 2827 -6750
rect 2861 -6784 2925 -6750
rect 2959 -6784 3023 -6750
rect 3057 -6784 3121 -6750
rect 3155 -6784 3219 -6750
rect 3253 -6784 3317 -6750
rect 3351 -6784 3415 -6750
rect 3449 -6784 3513 -6750
rect 3547 -6784 3611 -6750
rect 3645 -6784 3709 -6750
rect 3743 -6784 3807 -6750
rect 3841 -6784 3905 -6750
rect 3939 -6784 3955 -6750
rect 2517 -6892 2533 -6858
rect 2567 -6892 2631 -6858
rect 2665 -6892 2729 -6858
rect 2763 -6892 2827 -6858
rect 2861 -6892 2925 -6858
rect 2959 -6892 3023 -6858
rect 3057 -6892 3121 -6858
rect 3155 -6892 3219 -6858
rect 3253 -6892 3317 -6858
rect 3351 -6892 3415 -6858
rect 3449 -6892 3513 -6858
rect 3547 -6892 3611 -6858
rect 3645 -6892 3709 -6858
rect 3743 -6892 3807 -6858
rect 3841 -6892 3905 -6858
rect 3939 -6892 3955 -6858
rect 2484 -6942 2518 -6926
rect 2484 -7334 2518 -7318
rect 2582 -6942 2616 -6926
rect 2582 -7334 2616 -7318
rect 2680 -6942 2714 -6926
rect 2680 -7334 2714 -7318
rect 2778 -6942 2812 -6926
rect 2778 -7334 2812 -7318
rect 2876 -6942 2910 -6926
rect 2876 -7334 2910 -7318
rect 2974 -6942 3008 -6926
rect 2974 -7334 3008 -7318
rect 3072 -6942 3106 -6926
rect 3072 -7334 3106 -7318
rect 3170 -6942 3204 -6926
rect 3170 -7334 3204 -7318
rect 3268 -6942 3302 -6926
rect 3268 -7334 3302 -7318
rect 3366 -6942 3400 -6926
rect 3366 -7334 3400 -7318
rect 3464 -6942 3498 -6926
rect 3464 -7334 3498 -7318
rect 3562 -6942 3596 -6926
rect 3562 -7334 3596 -7318
rect 3660 -6942 3694 -6926
rect 3660 -7334 3694 -7318
rect 3758 -6942 3792 -6926
rect 3758 -7334 3792 -7318
rect 3856 -6942 3890 -6926
rect 3856 -7334 3890 -7318
rect 3954 -6942 3988 -6926
rect 3954 -7334 3988 -7318
rect 2517 -7402 2533 -7368
rect 2567 -7402 2631 -7368
rect 2665 -7402 2729 -7368
rect 2763 -7402 2827 -7368
rect 2861 -7402 2925 -7368
rect 2959 -7402 3023 -7368
rect 3057 -7402 3121 -7368
rect 3155 -7402 3219 -7368
rect 3253 -7402 3317 -7368
rect 3351 -7402 3415 -7368
rect 3449 -7402 3513 -7368
rect 3547 -7402 3611 -7368
rect 3645 -7402 3709 -7368
rect 3743 -7402 3807 -7368
rect 3841 -7402 3905 -7368
rect 3939 -7402 3955 -7368
rect 2294 -7470 2404 -7408
rect 4102 -7408 4174 -6940
rect 4068 -7470 4174 -7408
rect 2294 -7504 2466 -7470
rect 4006 -7504 4174 -7470
rect 2294 -7570 4174 -7504
rect 2071 -7769 2105 -7743
rect 4363 -7769 4397 -7743
rect 2071 -7803 2131 -7769
rect 4337 -7803 4397 -7769
rect 4800 -7916 5340 -2570
rect 1422 -7950 1596 -7916
rect 2818 -7950 2914 -7916
rect 1422 -8012 1534 -7950
rect 1422 -8532 1500 -8012
rect 1388 -8568 1500 -8532
rect 2880 -8012 2914 -7950
rect 1646 -8052 1662 -8018
rect 1696 -8052 1758 -8018
rect 1792 -8052 1854 -8018
rect 1888 -8052 1950 -8018
rect 1984 -8052 2046 -8018
rect 2080 -8052 2142 -8018
rect 2176 -8052 2238 -8018
rect 2272 -8052 2334 -8018
rect 2368 -8052 2430 -8018
rect 2464 -8052 2526 -8018
rect 2560 -8052 2622 -8018
rect 2656 -8052 2718 -8018
rect 2752 -8052 2768 -8018
rect 1614 -8102 1648 -8086
rect 1614 -8494 1648 -8478
rect 1710 -8102 1744 -8086
rect 1710 -8494 1744 -8478
rect 1806 -8102 1840 -8086
rect 1806 -8494 1840 -8478
rect 1902 -8102 1936 -8086
rect 1902 -8494 1936 -8478
rect 1998 -8102 2032 -8086
rect 1998 -8494 2032 -8478
rect 2094 -8102 2128 -8086
rect 2094 -8494 2128 -8478
rect 2190 -8102 2224 -8086
rect 2190 -8494 2224 -8478
rect 2286 -8102 2320 -8086
rect 2286 -8494 2320 -8478
rect 2382 -8102 2416 -8086
rect 2382 -8494 2416 -8478
rect 2478 -8102 2512 -8086
rect 2478 -8494 2512 -8478
rect 2574 -8102 2608 -8086
rect 2574 -8494 2608 -8478
rect 2670 -8102 2704 -8086
rect 2670 -8494 2704 -8478
rect 2766 -8102 2800 -8086
rect 2766 -8494 2800 -8478
rect 1646 -8562 1662 -8528
rect 1696 -8562 1758 -8528
rect 1792 -8562 1854 -8528
rect 1888 -8562 1950 -8528
rect 1984 -8562 2046 -8528
rect 2080 -8562 2142 -8528
rect 2176 -8562 2238 -8528
rect 2272 -8562 2334 -8528
rect 2368 -8562 2430 -8528
rect 2464 -8562 2526 -8528
rect 2560 -8562 2622 -8528
rect 2656 -8562 2718 -8528
rect 2752 -8562 2768 -8528
rect 1388 -8594 1534 -8568
rect -1396 -8628 -1194 -8594
rect 1326 -8628 1534 -8594
rect -1396 -8630 1534 -8628
rect 2880 -8630 2914 -8568
rect -1396 -8664 1596 -8630
rect 2818 -8664 2914 -8630
rect 3396 -7950 3492 -7916
rect 4714 -7950 5340 -7916
rect 3396 -8012 3430 -7950
rect 4776 -8012 5340 -7950
rect 3542 -8052 3558 -8018
rect 3592 -8052 3654 -8018
rect 3688 -8052 3750 -8018
rect 3784 -8052 3846 -8018
rect 3880 -8052 3942 -8018
rect 3976 -8052 4038 -8018
rect 4072 -8052 4134 -8018
rect 4168 -8052 4230 -8018
rect 4264 -8052 4326 -8018
rect 4360 -8052 4422 -8018
rect 4456 -8052 4518 -8018
rect 4552 -8052 4614 -8018
rect 4648 -8052 4664 -8018
rect 3510 -8102 3544 -8086
rect 3510 -8494 3544 -8478
rect 3606 -8102 3640 -8086
rect 3606 -8494 3640 -8478
rect 3702 -8102 3736 -8086
rect 3702 -8494 3736 -8478
rect 3798 -8102 3832 -8086
rect 3798 -8494 3832 -8478
rect 3894 -8102 3928 -8086
rect 3894 -8494 3928 -8478
rect 3990 -8102 4024 -8086
rect 3990 -8494 4024 -8478
rect 4086 -8102 4120 -8086
rect 4086 -8494 4120 -8478
rect 4182 -8102 4216 -8086
rect 4182 -8494 4216 -8478
rect 4278 -8102 4312 -8086
rect 4278 -8494 4312 -8478
rect 4374 -8102 4408 -8086
rect 4374 -8494 4408 -8478
rect 4470 -8102 4504 -8086
rect 4470 -8494 4504 -8478
rect 4566 -8102 4600 -8086
rect 4566 -8494 4600 -8478
rect 4662 -8102 4696 -8086
rect 4662 -8494 4696 -8478
rect 3542 -8562 3558 -8528
rect 3592 -8562 3654 -8528
rect 3688 -8562 3750 -8528
rect 3784 -8562 3846 -8528
rect 3880 -8562 3942 -8528
rect 3976 -8562 4038 -8528
rect 4072 -8562 4134 -8528
rect 4168 -8562 4230 -8528
rect 4264 -8562 4326 -8528
rect 4360 -8562 4422 -8528
rect 4456 -8562 4518 -8528
rect 4552 -8562 4614 -8528
rect 4648 -8562 4664 -8528
rect 3396 -8630 3430 -8568
rect 4810 -8568 5340 -8012
rect 4776 -8630 5340 -8568
rect 3396 -8660 3492 -8630
rect -1396 -8682 2914 -8664
rect -1396 -8716 -1214 -8682
rect 1256 -8716 2914 -8682
rect -1396 -8778 -1256 -8716
rect -1396 -11188 -1310 -8778
rect -1276 -11188 -1256 -8778
rect 1318 -8736 2914 -8716
rect 3300 -8664 3492 -8660
rect 4714 -8664 5340 -8630
rect 3300 -8730 5340 -8664
rect 3300 -8736 5390 -8730
rect 1318 -8770 1596 -8736
rect 3214 -8770 3492 -8736
rect 5110 -8770 5442 -8736
rect 5992 -8770 6088 -8736
rect 1318 -8778 1534 -8770
rect -1164 -8818 -1148 -8784
rect -1114 -8818 -1098 -8784
rect -972 -8818 -956 -8784
rect -922 -8818 -906 -8784
rect -780 -8818 -764 -8784
rect -730 -8818 -714 -8784
rect -588 -8818 -572 -8784
rect -538 -8818 -522 -8784
rect -396 -8818 -380 -8784
rect -346 -8818 -330 -8784
rect -204 -8818 -188 -8784
rect -154 -8818 -138 -8784
rect -12 -8818 4 -8784
rect 38 -8818 54 -8784
rect 180 -8818 196 -8784
rect 230 -8818 246 -8784
rect 372 -8818 388 -8784
rect 422 -8818 438 -8784
rect 564 -8818 580 -8784
rect 614 -8818 630 -8784
rect 756 -8818 772 -8784
rect 806 -8818 822 -8784
rect 948 -8818 964 -8784
rect 998 -8818 1014 -8784
rect 1140 -8818 1156 -8784
rect 1190 -8818 1206 -8784
rect -1196 -8868 -1162 -8852
rect -1196 -9260 -1162 -9244
rect -1100 -8868 -1066 -8852
rect -1100 -9260 -1066 -9244
rect -1004 -8868 -970 -8852
rect -1004 -9260 -970 -9244
rect -908 -8868 -874 -8852
rect -908 -9260 -874 -9244
rect -812 -8868 -778 -8852
rect -812 -9260 -778 -9244
rect -716 -8868 -682 -8852
rect -716 -9260 -682 -9244
rect -620 -8868 -586 -8852
rect -620 -9260 -586 -9244
rect -524 -8868 -490 -8852
rect -524 -9260 -490 -9244
rect -428 -8868 -394 -8852
rect -428 -9260 -394 -9244
rect -332 -8868 -298 -8852
rect -332 -9260 -298 -9244
rect -236 -8868 -202 -8852
rect -236 -9260 -202 -9244
rect -140 -8868 -106 -8852
rect -140 -9260 -106 -9244
rect -44 -8868 -10 -8852
rect -44 -9260 -10 -9244
rect 52 -8868 86 -8852
rect 52 -9260 86 -9244
rect 148 -8868 182 -8852
rect 148 -9260 182 -9244
rect 244 -8868 278 -8852
rect 244 -9260 278 -9244
rect 340 -8868 374 -8852
rect 340 -9260 374 -9244
rect 436 -8868 470 -8852
rect 436 -9260 470 -9244
rect 532 -8868 566 -8852
rect 532 -9260 566 -9244
rect 628 -8868 662 -8852
rect 628 -9260 662 -9244
rect 724 -8868 758 -8852
rect 724 -9260 758 -9244
rect 820 -8868 854 -8852
rect 820 -9260 854 -9244
rect 916 -8868 950 -8852
rect 916 -9260 950 -9244
rect 1012 -8868 1046 -8852
rect 1012 -9260 1046 -9244
rect 1108 -8868 1142 -8852
rect 1108 -9260 1142 -9244
rect 1204 -8868 1238 -8852
rect 1204 -9260 1238 -9244
rect 1352 -8832 1534 -8778
rect 1352 -9140 1500 -8832
rect -1068 -9328 -1052 -9294
rect -1018 -9328 -1002 -9294
rect -876 -9328 -860 -9294
rect -826 -9328 -810 -9294
rect -684 -9328 -668 -9294
rect -634 -9328 -618 -9294
rect -492 -9328 -476 -9294
rect -442 -9328 -426 -9294
rect -300 -9328 -284 -9294
rect -250 -9328 -234 -9294
rect -108 -9328 -92 -9294
rect -58 -9328 -42 -9294
rect 84 -9328 100 -9294
rect 134 -9328 150 -9294
rect 276 -9328 292 -9294
rect 326 -9328 342 -9294
rect 468 -9328 484 -9294
rect 518 -9328 534 -9294
rect 660 -9328 676 -9294
rect 710 -9328 726 -9294
rect 852 -9328 868 -9294
rect 902 -9328 918 -9294
rect 1044 -9328 1060 -9294
rect 1094 -9328 1110 -9294
rect 1474 -9320 1500 -9140
rect -1068 -9436 -1052 -9402
rect -1018 -9436 -1002 -9402
rect -876 -9436 -860 -9402
rect -826 -9436 -810 -9402
rect -684 -9436 -668 -9402
rect -634 -9436 -618 -9402
rect -492 -9436 -476 -9402
rect -442 -9436 -426 -9402
rect -300 -9436 -284 -9402
rect -250 -9436 -234 -9402
rect -108 -9436 -92 -9402
rect -58 -9436 -42 -9402
rect 84 -9436 100 -9402
rect 134 -9436 150 -9402
rect 276 -9436 292 -9402
rect 326 -9436 342 -9402
rect 468 -9436 484 -9402
rect 518 -9436 534 -9402
rect 660 -9436 676 -9402
rect 710 -9436 726 -9402
rect 852 -9436 868 -9402
rect 902 -9436 918 -9402
rect 1044 -9436 1060 -9402
rect 1094 -9436 1110 -9402
rect -1196 -9486 -1162 -9470
rect -1196 -9878 -1162 -9862
rect -1100 -9486 -1066 -9470
rect -1100 -9878 -1066 -9862
rect -1004 -9486 -970 -9470
rect -1004 -9878 -970 -9862
rect -908 -9486 -874 -9470
rect -908 -9878 -874 -9862
rect -812 -9486 -778 -9470
rect -812 -9878 -778 -9862
rect -716 -9486 -682 -9470
rect -716 -9878 -682 -9862
rect -620 -9486 -586 -9470
rect -620 -9878 -586 -9862
rect -524 -9486 -490 -9470
rect -524 -9878 -490 -9862
rect -428 -9486 -394 -9470
rect -428 -9878 -394 -9862
rect -332 -9486 -298 -9470
rect -332 -9878 -298 -9862
rect -236 -9486 -202 -9470
rect -236 -9878 -202 -9862
rect -140 -9486 -106 -9470
rect -140 -9878 -106 -9862
rect -44 -9486 -10 -9470
rect -44 -9878 -10 -9862
rect 52 -9486 86 -9470
rect 52 -9878 86 -9862
rect 148 -9486 182 -9470
rect 148 -9878 182 -9862
rect 244 -9486 278 -9470
rect 244 -9878 278 -9862
rect 340 -9486 374 -9470
rect 340 -9878 374 -9862
rect 436 -9486 470 -9470
rect 436 -9878 470 -9862
rect 532 -9486 566 -9470
rect 532 -9878 566 -9862
rect 628 -9486 662 -9470
rect 628 -9878 662 -9862
rect 724 -9486 758 -9470
rect 724 -9878 758 -9862
rect 820 -9486 854 -9470
rect 820 -9878 854 -9862
rect 916 -9486 950 -9470
rect 916 -9878 950 -9862
rect 1012 -9486 1046 -9470
rect 1012 -9878 1046 -9862
rect 1108 -9486 1142 -9470
rect 1108 -9878 1142 -9862
rect 1204 -9486 1238 -9470
rect 1204 -9878 1238 -9862
rect -1164 -9946 -1148 -9912
rect -1114 -9946 -1098 -9912
rect -972 -9946 -956 -9912
rect -922 -9946 -906 -9912
rect -780 -9946 -764 -9912
rect -730 -9946 -714 -9912
rect -588 -9946 -572 -9912
rect -538 -9946 -522 -9912
rect -396 -9946 -380 -9912
rect -346 -9946 -330 -9912
rect -204 -9946 -188 -9912
rect -154 -9946 -138 -9912
rect -12 -9946 4 -9912
rect 38 -9946 54 -9912
rect 180 -9946 196 -9912
rect 230 -9946 246 -9912
rect 372 -9946 388 -9912
rect 422 -9946 438 -9912
rect 564 -9946 580 -9912
rect 614 -9946 630 -9912
rect 756 -9946 772 -9912
rect 806 -9946 822 -9912
rect 948 -9946 964 -9912
rect 998 -9946 1014 -9912
rect 1140 -9946 1156 -9912
rect 1190 -9946 1206 -9912
rect -1164 -10054 -1148 -10020
rect -1114 -10054 -1098 -10020
rect -972 -10054 -956 -10020
rect -922 -10054 -906 -10020
rect -780 -10054 -764 -10020
rect -730 -10054 -714 -10020
rect -588 -10054 -572 -10020
rect -538 -10054 -522 -10020
rect -396 -10054 -380 -10020
rect -346 -10054 -330 -10020
rect -204 -10054 -188 -10020
rect -154 -10054 -138 -10020
rect -12 -10054 4 -10020
rect 38 -10054 54 -10020
rect 180 -10054 196 -10020
rect 230 -10054 246 -10020
rect 372 -10054 388 -10020
rect 422 -10054 438 -10020
rect 564 -10054 580 -10020
rect 614 -10054 630 -10020
rect 756 -10054 772 -10020
rect 806 -10054 822 -10020
rect 948 -10054 964 -10020
rect 998 -10054 1014 -10020
rect 1140 -10054 1156 -10020
rect 1190 -10054 1206 -10020
rect -1196 -10104 -1162 -10088
rect -1196 -10496 -1162 -10480
rect -1100 -10104 -1066 -10088
rect -1100 -10496 -1066 -10480
rect -1004 -10104 -970 -10088
rect -1004 -10496 -970 -10480
rect -908 -10104 -874 -10088
rect -908 -10496 -874 -10480
rect -812 -10104 -778 -10088
rect -812 -10496 -778 -10480
rect -716 -10104 -682 -10088
rect -716 -10496 -682 -10480
rect -620 -10104 -586 -10088
rect -620 -10496 -586 -10480
rect -524 -10104 -490 -10088
rect -524 -10496 -490 -10480
rect -428 -10104 -394 -10088
rect -428 -10496 -394 -10480
rect -332 -10104 -298 -10088
rect -332 -10496 -298 -10480
rect -236 -10104 -202 -10088
rect -236 -10496 -202 -10480
rect -140 -10104 -106 -10088
rect -140 -10496 -106 -10480
rect -44 -10104 -10 -10088
rect -44 -10496 -10 -10480
rect 52 -10104 86 -10088
rect 52 -10496 86 -10480
rect 148 -10104 182 -10088
rect 148 -10496 182 -10480
rect 244 -10104 278 -10088
rect 244 -10496 278 -10480
rect 340 -10104 374 -10088
rect 340 -10496 374 -10480
rect 436 -10104 470 -10088
rect 436 -10496 470 -10480
rect 532 -10104 566 -10088
rect 532 -10496 566 -10480
rect 628 -10104 662 -10088
rect 628 -10496 662 -10480
rect 724 -10104 758 -10088
rect 724 -10496 758 -10480
rect 820 -10104 854 -10088
rect 820 -10496 854 -10480
rect 916 -10104 950 -10088
rect 916 -10496 950 -10480
rect 1012 -10104 1046 -10088
rect 1012 -10496 1046 -10480
rect 1108 -10104 1142 -10088
rect 1108 -10496 1142 -10480
rect 1204 -10104 1238 -10088
rect 1204 -10496 1238 -10480
rect -1068 -10564 -1052 -10530
rect -1018 -10564 -1002 -10530
rect -876 -10564 -860 -10530
rect -826 -10564 -810 -10530
rect -684 -10564 -668 -10530
rect -634 -10564 -618 -10530
rect -492 -10564 -476 -10530
rect -442 -10564 -426 -10530
rect -300 -10564 -284 -10530
rect -250 -10564 -234 -10530
rect -108 -10564 -92 -10530
rect -58 -10564 -42 -10530
rect 84 -10564 100 -10530
rect 134 -10564 150 -10530
rect 276 -10564 292 -10530
rect 326 -10564 342 -10530
rect 468 -10564 484 -10530
rect 518 -10564 534 -10530
rect 660 -10564 676 -10530
rect 710 -10564 726 -10530
rect 852 -10564 868 -10530
rect 902 -10564 918 -10530
rect 1044 -10564 1060 -10530
rect 1094 -10564 1110 -10530
rect -1068 -10672 -1052 -10638
rect -1018 -10672 -1002 -10638
rect -876 -10672 -860 -10638
rect -826 -10672 -810 -10638
rect -684 -10672 -668 -10638
rect -634 -10672 -618 -10638
rect -492 -10672 -476 -10638
rect -442 -10672 -426 -10638
rect -300 -10672 -284 -10638
rect -250 -10672 -234 -10638
rect -108 -10672 -92 -10638
rect -58 -10672 -42 -10638
rect 84 -10672 100 -10638
rect 134 -10672 150 -10638
rect 276 -10672 292 -10638
rect 326 -10672 342 -10638
rect 468 -10672 484 -10638
rect 518 -10672 534 -10638
rect 660 -10672 676 -10638
rect 710 -10672 726 -10638
rect 852 -10672 868 -10638
rect 902 -10672 918 -10638
rect 1044 -10672 1060 -10638
rect 1094 -10672 1110 -10638
rect -1196 -10722 -1162 -10706
rect -1196 -11114 -1162 -11098
rect -1100 -10722 -1066 -10706
rect -1100 -11114 -1066 -11098
rect -1004 -10722 -970 -10706
rect -1004 -11114 -970 -11098
rect -908 -10722 -874 -10706
rect -908 -11114 -874 -11098
rect -812 -10722 -778 -10706
rect -812 -11114 -778 -11098
rect -716 -10722 -682 -10706
rect -716 -11114 -682 -11098
rect -620 -10722 -586 -10706
rect -620 -11114 -586 -11098
rect -524 -10722 -490 -10706
rect -524 -11114 -490 -11098
rect -428 -10722 -394 -10706
rect -428 -11114 -394 -11098
rect -332 -10722 -298 -10706
rect -332 -11114 -298 -11098
rect -236 -10722 -202 -10706
rect -236 -11114 -202 -11098
rect -140 -10722 -106 -10706
rect -140 -11114 -106 -11098
rect -44 -10722 -10 -10706
rect -44 -11114 -10 -11098
rect 52 -10722 86 -10706
rect 52 -11114 86 -11098
rect 148 -10722 182 -10706
rect 148 -11114 182 -11098
rect 244 -10722 278 -10706
rect 244 -11114 278 -11098
rect 340 -10722 374 -10706
rect 340 -11114 374 -11098
rect 436 -10722 470 -10706
rect 436 -11114 470 -11098
rect 532 -10722 566 -10706
rect 532 -11114 566 -11098
rect 628 -10722 662 -10706
rect 628 -11114 662 -11098
rect 724 -10722 758 -10706
rect 724 -11114 758 -11098
rect 820 -10722 854 -10706
rect 820 -11114 854 -11098
rect 916 -10722 950 -10706
rect 916 -11114 950 -11098
rect 1012 -10722 1046 -10706
rect 1012 -11114 1046 -11098
rect 1108 -10722 1142 -10706
rect 1108 -11114 1142 -11098
rect 1204 -10722 1238 -10706
rect 1204 -11114 1238 -11098
rect -1164 -11182 -1148 -11148
rect -1114 -11182 -1098 -11148
rect -972 -11182 -956 -11148
rect -922 -11182 -906 -11148
rect -780 -11182 -764 -11148
rect -730 -11182 -714 -11148
rect -588 -11182 -572 -11148
rect -538 -11182 -522 -11148
rect -396 -11182 -380 -11148
rect -346 -11182 -330 -11148
rect -204 -11182 -188 -11148
rect -154 -11182 -138 -11148
rect -12 -11182 4 -11148
rect 38 -11182 54 -11148
rect 180 -11182 196 -11148
rect 230 -11182 246 -11148
rect 372 -11182 388 -11148
rect 422 -11182 438 -11148
rect 564 -11182 580 -11148
rect 614 -11182 630 -11148
rect 756 -11182 772 -11148
rect 806 -11182 822 -11148
rect 948 -11182 964 -11148
rect 998 -11182 1014 -11148
rect 1140 -11182 1156 -11148
rect 1190 -11182 1206 -11148
rect -1396 -11250 -1256 -11188
rect 1352 -9388 1500 -9320
rect 3276 -8832 3430 -8770
rect 1660 -8872 1676 -8838
rect 1844 -8872 1860 -8838
rect 1918 -8872 1934 -8838
rect 2102 -8872 2118 -8838
rect 2176 -8872 2192 -8838
rect 2360 -8872 2376 -8838
rect 2434 -8872 2450 -8838
rect 2618 -8872 2634 -8838
rect 2692 -8872 2708 -8838
rect 2876 -8872 2892 -8838
rect 2950 -8872 2966 -8838
rect 3134 -8872 3150 -8838
rect 1614 -8922 1648 -8906
rect 1614 -9314 1648 -9298
rect 1872 -8922 1906 -8906
rect 1872 -9314 1906 -9298
rect 2130 -8922 2164 -8906
rect 2130 -9314 2164 -9298
rect 2388 -8922 2422 -8906
rect 2388 -9314 2422 -9298
rect 2646 -8922 2680 -8906
rect 2646 -9314 2680 -9298
rect 2904 -8922 2938 -8906
rect 2904 -9314 2938 -9298
rect 3162 -8922 3196 -8906
rect 3162 -9314 3196 -9298
rect 1660 -9382 1676 -9348
rect 1844 -9382 1860 -9348
rect 1918 -9382 1934 -9348
rect 2102 -9382 2118 -9348
rect 2176 -9382 2192 -9348
rect 2360 -9382 2376 -9348
rect 2434 -9382 2450 -9348
rect 2618 -9382 2634 -9348
rect 2692 -9382 2708 -9348
rect 2876 -9382 2892 -9348
rect 2950 -9382 2966 -9348
rect 3134 -9382 3150 -9348
rect 1352 -9450 1534 -9388
rect 3310 -9388 3396 -8832
rect 5172 -8832 5380 -8770
rect 3556 -8872 3572 -8838
rect 3740 -8872 3756 -8838
rect 3814 -8872 3830 -8838
rect 3998 -8872 4014 -8838
rect 4072 -8872 4088 -8838
rect 4256 -8872 4272 -8838
rect 4330 -8872 4346 -8838
rect 4514 -8872 4530 -8838
rect 4588 -8872 4604 -8838
rect 4772 -8872 4788 -8838
rect 4846 -8872 4862 -8838
rect 5030 -8872 5046 -8838
rect 3510 -8922 3544 -8906
rect 3510 -9314 3544 -9298
rect 3768 -8922 3802 -8906
rect 3768 -9314 3802 -9298
rect 4026 -8922 4060 -8906
rect 4026 -9314 4060 -9298
rect 4284 -8922 4318 -8906
rect 4284 -9314 4318 -9298
rect 4542 -8922 4576 -8906
rect 4542 -9314 4576 -9298
rect 4800 -8922 4834 -8906
rect 4800 -9314 4834 -9298
rect 5058 -8922 5092 -8906
rect 5058 -9314 5092 -9298
rect 3556 -9382 3572 -9348
rect 3740 -9382 3756 -9348
rect 3814 -9382 3830 -9348
rect 3998 -9382 4014 -9348
rect 4072 -9382 4088 -9348
rect 4256 -9382 4272 -9348
rect 4330 -9382 4346 -9348
rect 4514 -9382 4530 -9348
rect 4588 -9382 4604 -9348
rect 4772 -9382 4788 -9348
rect 4846 -9382 4862 -9348
rect 5030 -9382 5046 -9348
rect 3276 -9450 3430 -9388
rect 5206 -9388 5346 -8832
rect 6054 -8832 6088 -8770
rect 5588 -8872 5604 -8838
rect 5638 -8872 5654 -8838
rect 5780 -8872 5796 -8838
rect 5830 -8872 5846 -8838
rect 5460 -8922 5494 -8906
rect 5460 -9314 5494 -9298
rect 5556 -8922 5590 -8906
rect 5556 -9314 5590 -9298
rect 5652 -8922 5686 -8906
rect 5652 -9314 5686 -9298
rect 5748 -8922 5782 -8906
rect 5748 -9314 5782 -9298
rect 5844 -8922 5878 -8906
rect 5844 -9314 5878 -9298
rect 5940 -8922 5974 -8906
rect 5974 -9298 6054 -9150
rect 5940 -9314 6054 -9298
rect 5970 -9320 6054 -9314
rect 5492 -9382 5508 -9348
rect 5542 -9382 5558 -9348
rect 5684 -9382 5700 -9348
rect 5734 -9382 5750 -9348
rect 5876 -9382 5892 -9348
rect 5926 -9382 5942 -9348
rect 5172 -9450 5380 -9388
rect 5980 -9388 6054 -9320
rect 5980 -9450 6088 -9388
rect 1352 -9484 1596 -9450
rect 3214 -9484 3492 -9450
rect 5110 -9484 5442 -9450
rect 5992 -9470 6088 -9450
rect 5992 -9484 6090 -9470
rect 1352 -9730 6090 -9484
rect 1352 -9764 1582 -9730
rect 5884 -9740 6090 -9730
rect 5884 -9764 5980 -9740
rect 1352 -9853 1520 -9764
rect 1352 -10991 1486 -9853
rect 1693 -9884 1709 -9850
rect 2077 -9884 2093 -9850
rect 2160 -9930 2540 -9764
rect 2613 -9884 2629 -9850
rect 2997 -9884 3013 -9850
rect 3070 -9930 3450 -9764
rect 3533 -9884 3549 -9850
rect 3917 -9884 3933 -9850
rect 4000 -9930 4380 -9764
rect 4453 -9884 4469 -9850
rect 4837 -9884 4853 -9850
rect 4910 -9930 5310 -9764
rect 5373 -9884 5389 -9850
rect 5757 -9884 5773 -9850
rect 5840 -9853 5980 -9764
rect 5840 -9930 5946 -9853
rect 1608 -9946 1642 -9930
rect 1608 -10914 1642 -10898
rect 2144 -9946 2562 -9930
rect 2178 -10898 2528 -9946
rect 2144 -10914 2562 -10898
rect 3064 -9946 3482 -9930
rect 3098 -10898 3448 -9946
rect 3064 -10914 3482 -10898
rect 3984 -9946 4402 -9930
rect 4018 -10898 4368 -9946
rect 3984 -10914 4402 -10898
rect 4904 -9946 5322 -9930
rect 4938 -10898 5288 -9946
rect 4904 -10914 5322 -10898
rect 5824 -9946 5946 -9930
rect 5858 -10898 5946 -9946
rect 5824 -10914 5946 -10898
rect 1352 -11080 1520 -10991
rect 1693 -10994 1709 -10960
rect 2077 -10994 2093 -10960
rect 2160 -11080 2540 -10914
rect 2613 -10994 2629 -10960
rect 2997 -10994 3013 -10960
rect 3070 -11080 3450 -10914
rect 3533 -10994 3549 -10960
rect 3917 -10994 3933 -10960
rect 4000 -11080 4380 -10914
rect 4453 -10994 4469 -10960
rect 4837 -10994 4853 -10960
rect 4910 -11080 5310 -10914
rect 5373 -10994 5389 -10960
rect 5757 -10994 5773 -10960
rect 5840 -10991 5946 -10914
rect 6216 -10062 6312 -10028
rect 6640 -10062 6736 -10028
rect 6216 -10124 6250 -10062
rect 6702 -10124 6736 -10062
rect 6376 -10164 6392 -10130
rect 6560 -10164 6576 -10130
rect 6620 -10207 6670 -10200
rect 6330 -10223 6364 -10207
rect 6330 -10315 6364 -10299
rect 6588 -10223 6670 -10207
rect 6622 -10299 6670 -10223
rect 6588 -10315 6670 -10299
rect 6620 -10320 6670 -10315
rect 6376 -10392 6392 -10358
rect 6560 -10392 6576 -10358
rect 6216 -10460 6250 -10398
rect 6702 -10460 6736 -10398
rect 6216 -10494 6312 -10460
rect 6640 -10494 6736 -10460
rect 6216 -10600 6312 -10596
rect 5980 -10630 6312 -10600
rect 6640 -10630 6736 -10596
rect 5980 -10692 6250 -10630
rect 5980 -10948 6216 -10692
rect 6702 -10692 6736 -10630
rect 6376 -10732 6392 -10698
rect 6560 -10732 6576 -10698
rect 6610 -10766 6702 -10760
rect 6330 -10782 6364 -10766
rect 6330 -10874 6364 -10858
rect 6588 -10782 6702 -10766
rect 6622 -10858 6702 -10782
rect 6588 -10874 6702 -10858
rect 6610 -10880 6702 -10874
rect 6376 -10942 6392 -10908
rect 6560 -10942 6576 -10908
rect 5980 -10991 6250 -10948
rect 5840 -11010 6250 -10991
rect 6702 -11010 6736 -10948
rect 5840 -11040 6312 -11010
rect 5840 -11080 5980 -11040
rect 6216 -11044 6312 -11040
rect 6640 -11044 6736 -11010
rect 1352 -11114 1609 -11080
rect 5857 -11114 5980 -11080
rect 1352 -11188 5970 -11114
rect 1318 -11250 5970 -11188
rect -1396 -11284 -1214 -11250
rect 1256 -11280 5970 -11250
rect 1256 -11284 1352 -11280
rect -1396 -11290 -1256 -11284
<< viali >>
rect -1127 2592 -1093 2626
rect -1029 2592 -995 2626
rect -931 2592 -897 2626
rect -833 2592 -799 2626
rect -735 2592 -701 2626
rect -637 2592 -603 2626
rect -539 2592 -505 2626
rect -441 2592 -407 2626
rect -343 2592 -309 2626
rect -245 2592 -211 2626
rect -147 2592 -113 2626
rect -49 2592 -15 2626
rect 49 2592 83 2626
rect 147 2592 181 2626
rect 245 2592 279 2626
rect -1176 2157 -1142 2533
rect -1078 2157 -1044 2533
rect -980 2157 -946 2533
rect -882 2157 -848 2533
rect -784 2157 -750 2533
rect -686 2157 -652 2533
rect -588 2157 -554 2533
rect -490 2157 -456 2533
rect -392 2157 -358 2533
rect -294 2157 -260 2533
rect -196 2157 -162 2533
rect -98 2157 -64 2533
rect 0 2157 34 2533
rect 98 2157 132 2533
rect 196 2157 230 2533
rect 294 2157 328 2533
rect -1127 2064 -1093 2098
rect -1029 2064 -995 2098
rect -931 2064 -897 2098
rect -833 2064 -799 2098
rect -735 2064 -701 2098
rect -637 2064 -603 2098
rect -539 2064 -505 2098
rect -441 2064 -407 2098
rect -343 2064 -309 2098
rect -245 2064 -211 2098
rect -147 2064 -113 2098
rect -49 2064 -15 2098
rect 49 2064 83 2098
rect 147 2064 181 2098
rect 245 2064 279 2098
rect -1127 1956 -1093 1990
rect -1029 1956 -995 1990
rect -931 1956 -897 1990
rect -833 1956 -799 1990
rect -735 1956 -701 1990
rect -637 1956 -603 1990
rect -539 1956 -505 1990
rect -441 1956 -407 1990
rect -343 1956 -309 1990
rect -245 1956 -211 1990
rect -147 1956 -113 1990
rect -49 1956 -15 1990
rect 49 1956 83 1990
rect 147 1956 181 1990
rect 245 1956 279 1990
rect -1176 1521 -1142 1897
rect -1078 1521 -1044 1897
rect -980 1521 -946 1897
rect -882 1521 -848 1897
rect -784 1521 -750 1897
rect -686 1521 -652 1897
rect -588 1521 -554 1897
rect -490 1521 -456 1897
rect -392 1521 -358 1897
rect -294 1521 -260 1897
rect -196 1521 -162 1897
rect -98 1521 -64 1897
rect 0 1521 34 1897
rect 98 1521 132 1897
rect 196 1521 230 1897
rect 294 1521 328 1897
rect -1127 1428 -1093 1462
rect -1029 1428 -995 1462
rect -931 1428 -897 1462
rect -833 1428 -799 1462
rect -735 1428 -701 1462
rect -637 1428 -603 1462
rect -539 1428 -505 1462
rect -441 1428 -407 1462
rect -343 1428 -309 1462
rect -245 1428 -211 1462
rect -147 1428 -113 1462
rect -49 1428 -15 1462
rect 49 1428 83 1462
rect 147 1428 181 1462
rect 245 1428 279 1462
rect 671 2592 705 2626
rect 769 2592 803 2626
rect 867 2592 901 2626
rect 965 2592 999 2626
rect 1063 2592 1097 2626
rect 1161 2592 1195 2626
rect 1259 2592 1293 2626
rect 1357 2592 1391 2626
rect 1455 2592 1489 2626
rect 1553 2592 1587 2626
rect 1651 2592 1685 2626
rect 1749 2592 1783 2626
rect 1847 2592 1881 2626
rect 1945 2592 1979 2626
rect 2043 2592 2077 2626
rect 622 2157 656 2533
rect 720 2157 754 2533
rect 818 2157 852 2533
rect 916 2157 950 2533
rect 1014 2157 1048 2533
rect 1112 2157 1146 2533
rect 1210 2157 1244 2533
rect 1308 2157 1342 2533
rect 1406 2157 1440 2533
rect 1504 2157 1538 2533
rect 1602 2157 1636 2533
rect 1700 2157 1734 2533
rect 1798 2157 1832 2533
rect 1896 2157 1930 2533
rect 1994 2157 2028 2533
rect 2092 2157 2126 2533
rect 671 2064 705 2098
rect 769 2064 803 2098
rect 867 2064 901 2098
rect 965 2064 999 2098
rect 1063 2064 1097 2098
rect 1161 2064 1195 2098
rect 1259 2064 1293 2098
rect 1357 2064 1391 2098
rect 1455 2064 1489 2098
rect 1553 2064 1587 2098
rect 1651 2064 1685 2098
rect 1749 2064 1783 2098
rect 1847 2064 1881 2098
rect 1945 2064 1979 2098
rect 2043 2064 2077 2098
rect 671 1956 705 1990
rect 769 1956 803 1990
rect 867 1956 901 1990
rect 965 1956 999 1990
rect 1063 1956 1097 1990
rect 1161 1956 1195 1990
rect 1259 1956 1293 1990
rect 1357 1956 1391 1990
rect 1455 1956 1489 1990
rect 1553 1956 1587 1990
rect 1651 1956 1685 1990
rect 1749 1956 1783 1990
rect 1847 1956 1881 1990
rect 1945 1956 1979 1990
rect 2043 1956 2077 1990
rect 622 1521 656 1897
rect 720 1521 754 1897
rect 818 1521 852 1897
rect 916 1521 950 1897
rect 1014 1521 1048 1897
rect 1112 1521 1146 1897
rect 1210 1521 1244 1897
rect 1308 1521 1342 1897
rect 1406 1521 1440 1897
rect 1504 1521 1538 1897
rect 1602 1521 1636 1897
rect 1700 1521 1734 1897
rect 1798 1521 1832 1897
rect 1896 1521 1930 1897
rect 1994 1521 2028 1897
rect 2092 1521 2126 1897
rect 2214 1510 2240 2070
rect 2240 1980 2344 2070
rect 2240 1510 2310 1980
rect 2310 1510 2344 1980
rect 2486 1940 2554 1974
rect 2644 1940 2712 1974
rect 2802 1940 2870 1974
rect 2960 1940 3028 1974
rect 3118 1940 3186 1974
rect 3276 1940 3344 1974
rect 3434 1940 3502 1974
rect 3592 1940 3660 1974
rect 3750 1940 3818 1974
rect 3908 1940 3976 1974
rect 671 1428 705 1462
rect 769 1428 803 1462
rect 867 1428 901 1462
rect 965 1428 999 1462
rect 1063 1428 1097 1462
rect 1161 1428 1195 1462
rect 1259 1428 1293 1462
rect 1357 1428 1391 1462
rect 1455 1428 1489 1462
rect 1553 1428 1587 1462
rect 1651 1428 1685 1462
rect 1749 1428 1783 1462
rect 1847 1428 1881 1462
rect 1945 1428 1979 1462
rect 2043 1428 2077 1462
rect 2424 1505 2458 1881
rect 2582 1505 2616 1881
rect 2740 1505 2774 1881
rect 2898 1505 2932 1881
rect 3056 1505 3090 1881
rect 3214 1505 3248 1881
rect 3372 1505 3406 1881
rect 3530 1505 3564 1881
rect 3688 1505 3722 1881
rect 3846 1505 3880 1881
rect 4004 1505 4038 1881
rect 2486 1412 2554 1446
rect 2644 1412 2712 1446
rect 2802 1412 2870 1446
rect 2960 1412 3028 1446
rect 3118 1412 3186 1446
rect 3276 1412 3344 1446
rect 3434 1412 3502 1446
rect 3592 1412 3660 1446
rect 3750 1412 3818 1446
rect 3908 1412 3976 1446
rect -1127 1116 -1093 1150
rect -1030 1116 -996 1150
rect -931 1116 -897 1150
rect -834 1116 -800 1150
rect -735 1116 -701 1150
rect -638 1116 -604 1150
rect -539 1116 -505 1150
rect -442 1116 -408 1150
rect -343 1116 -309 1150
rect -246 1116 -212 1150
rect -147 1116 -113 1150
rect -50 1116 -16 1150
rect 49 1116 83 1150
rect 146 1116 180 1150
rect 245 1116 279 1150
rect 342 1116 376 1150
rect 441 1116 475 1150
rect 538 1116 572 1150
rect 637 1116 671 1150
rect 734 1116 768 1150
rect 833 1116 867 1150
rect 930 1116 964 1150
rect 1029 1116 1063 1150
rect 1126 1116 1160 1150
rect 1225 1116 1259 1150
rect -1176 690 -1142 1066
rect -1078 690 -1044 1066
rect -980 690 -946 1066
rect -882 690 -848 1066
rect -784 690 -750 1066
rect -686 690 -652 1066
rect -588 690 -554 1066
rect -490 690 -456 1066
rect -392 690 -358 1066
rect -294 690 -260 1066
rect -196 690 -162 1066
rect -98 690 -64 1066
rect 0 690 34 1066
rect 98 690 132 1066
rect 196 690 230 1066
rect 294 690 328 1066
rect 392 690 426 1066
rect 490 690 524 1066
rect 588 690 622 1066
rect 686 690 720 1066
rect 784 690 818 1066
rect 882 690 916 1066
rect 980 690 1014 1066
rect 1078 690 1112 1066
rect 1176 690 1210 1066
rect 1274 690 1308 1066
rect -1128 606 -1094 640
rect -1029 606 -995 640
rect -932 606 -898 640
rect -833 606 -799 640
rect -736 606 -702 640
rect -637 606 -603 640
rect -540 606 -506 640
rect -441 606 -407 640
rect -344 606 -310 640
rect -245 606 -211 640
rect -148 606 -114 640
rect -49 606 -15 640
rect 48 606 82 640
rect 147 606 181 640
rect 244 606 278 640
rect 343 606 377 640
rect 440 606 474 640
rect 539 606 573 640
rect 636 606 670 640
rect 735 606 769 640
rect 832 606 866 640
rect 931 606 965 640
rect 1028 606 1062 640
rect 1127 606 1161 640
rect 1224 606 1258 640
rect -1127 498 -1093 532
rect -1029 498 -995 532
rect -931 498 -897 532
rect -833 498 -799 532
rect -735 498 -701 532
rect -637 498 -603 532
rect -539 498 -505 532
rect -441 498 -407 532
rect -343 498 -309 532
rect -245 498 -211 532
rect -147 498 -113 532
rect -49 498 -15 532
rect 49 498 83 532
rect 147 498 181 532
rect 245 498 279 532
rect 343 498 377 532
rect 441 498 475 532
rect 539 498 573 532
rect 637 498 671 532
rect 735 498 769 532
rect 833 498 867 532
rect 931 498 965 532
rect 1029 498 1063 532
rect 1127 498 1161 532
rect 1225 498 1259 532
rect -1176 72 -1142 448
rect -1078 72 -1044 448
rect -980 72 -946 448
rect -882 72 -848 448
rect -784 72 -750 448
rect -686 72 -652 448
rect -588 72 -554 448
rect -490 72 -456 448
rect -392 72 -358 448
rect -294 72 -260 448
rect -196 72 -162 448
rect -98 72 -64 448
rect 0 72 34 448
rect 98 72 132 448
rect 196 72 230 448
rect 294 72 328 448
rect 392 72 426 448
rect 490 72 524 448
rect 588 72 622 448
rect 686 72 720 448
rect 784 72 818 448
rect 882 72 916 448
rect 980 72 1014 448
rect 1078 72 1112 448
rect 1176 72 1210 448
rect 1274 72 1308 448
rect -1127 -12 -1093 22
rect -1029 -12 -995 22
rect -931 -12 -897 22
rect -833 -12 -799 22
rect -735 -12 -701 22
rect -637 -12 -603 22
rect -539 -12 -505 22
rect -441 -12 -407 22
rect -343 -12 -309 22
rect -245 -12 -211 22
rect -147 -12 -113 22
rect -49 -12 -15 22
rect 49 -12 83 22
rect 147 -12 181 22
rect 245 -12 279 22
rect 343 -12 377 22
rect 441 -12 475 22
rect 539 -12 573 22
rect 637 -12 671 22
rect 735 -12 769 22
rect 833 -12 867 22
rect 931 -12 965 22
rect 1029 -12 1063 22
rect 1127 -12 1161 22
rect 1225 -12 1259 22
rect -1127 -328 -1093 -294
rect -1030 -328 -996 -294
rect -931 -328 -897 -294
rect -834 -328 -800 -294
rect -735 -328 -701 -294
rect -638 -328 -604 -294
rect -539 -328 -505 -294
rect -442 -328 -408 -294
rect -343 -328 -309 -294
rect -246 -328 -212 -294
rect -147 -328 -113 -294
rect -50 -328 -16 -294
rect 49 -328 83 -294
rect 146 -328 180 -294
rect 245 -328 279 -294
rect 342 -328 376 -294
rect 441 -328 475 -294
rect 538 -328 572 -294
rect 637 -328 671 -294
rect 734 -328 768 -294
rect 833 -328 867 -294
rect 930 -328 964 -294
rect 1029 -328 1063 -294
rect 1126 -328 1160 -294
rect 1225 -328 1259 -294
rect -1176 -754 -1142 -378
rect -1078 -754 -1044 -378
rect -980 -754 -946 -378
rect -882 -754 -848 -378
rect -784 -754 -750 -378
rect -686 -754 -652 -378
rect -588 -754 -554 -378
rect -490 -754 -456 -378
rect -392 -754 -358 -378
rect -294 -754 -260 -378
rect -196 -754 -162 -378
rect -98 -754 -64 -378
rect 0 -754 34 -378
rect 98 -754 132 -378
rect 196 -754 230 -378
rect 294 -754 328 -378
rect 392 -754 426 -378
rect 490 -754 524 -378
rect 588 -754 622 -378
rect 686 -754 720 -378
rect 784 -754 818 -378
rect 882 -754 916 -378
rect 980 -754 1014 -378
rect 1078 -754 1112 -378
rect 1176 -754 1210 -378
rect 1274 -754 1308 -378
rect -1128 -838 -1094 -804
rect -1029 -838 -995 -804
rect -932 -838 -898 -804
rect -833 -838 -799 -804
rect -736 -838 -702 -804
rect -637 -838 -603 -804
rect -540 -838 -506 -804
rect -441 -838 -407 -804
rect -344 -838 -310 -804
rect -245 -838 -211 -804
rect -148 -838 -114 -804
rect -49 -838 -15 -804
rect 48 -838 82 -804
rect 147 -838 181 -804
rect 244 -838 278 -804
rect 343 -838 377 -804
rect 440 -838 474 -804
rect 539 -838 573 -804
rect 636 -838 670 -804
rect 735 -838 769 -804
rect 832 -838 866 -804
rect 931 -838 965 -804
rect 1028 -838 1062 -804
rect 1127 -838 1161 -804
rect 1224 -838 1258 -804
rect -1127 -946 -1093 -912
rect -1029 -946 -995 -912
rect -931 -946 -897 -912
rect -833 -946 -799 -912
rect -735 -946 -701 -912
rect -637 -946 -603 -912
rect -539 -946 -505 -912
rect -441 -946 -407 -912
rect -343 -946 -309 -912
rect -245 -946 -211 -912
rect -147 -946 -113 -912
rect -49 -946 -15 -912
rect 49 -946 83 -912
rect 147 -946 181 -912
rect 245 -946 279 -912
rect 343 -946 377 -912
rect 441 -946 475 -912
rect 539 -946 573 -912
rect 637 -946 671 -912
rect 735 -946 769 -912
rect 833 -946 867 -912
rect 931 -946 965 -912
rect 1029 -946 1063 -912
rect 1127 -946 1161 -912
rect 1225 -946 1259 -912
rect -1176 -1372 -1142 -996
rect -1078 -1372 -1044 -996
rect -980 -1372 -946 -996
rect -882 -1372 -848 -996
rect -784 -1372 -750 -996
rect -686 -1372 -652 -996
rect -588 -1372 -554 -996
rect -490 -1372 -456 -996
rect -392 -1372 -358 -996
rect -294 -1372 -260 -996
rect -196 -1372 -162 -996
rect -98 -1372 -64 -996
rect 0 -1372 34 -996
rect 98 -1372 132 -996
rect 196 -1372 230 -996
rect 294 -1372 328 -996
rect 392 -1372 426 -996
rect 490 -1372 524 -996
rect 588 -1372 622 -996
rect 686 -1372 720 -996
rect 784 -1372 818 -996
rect 882 -1372 916 -996
rect 980 -1372 1014 -996
rect 1078 -1372 1112 -996
rect 1176 -1372 1210 -996
rect 1274 -1372 1308 -996
rect -1127 -1456 -1093 -1422
rect -1029 -1456 -995 -1422
rect -931 -1456 -897 -1422
rect -833 -1456 -799 -1422
rect -735 -1456 -701 -1422
rect -637 -1456 -603 -1422
rect -539 -1456 -505 -1422
rect -441 -1456 -407 -1422
rect -343 -1456 -309 -1422
rect -245 -1456 -211 -1422
rect -147 -1456 -113 -1422
rect -49 -1456 -15 -1422
rect 49 -1456 83 -1422
rect 147 -1456 181 -1422
rect 245 -1456 279 -1422
rect 343 -1456 377 -1422
rect 441 -1456 475 -1422
rect 539 -1456 573 -1422
rect 637 -1456 671 -1422
rect 735 -1456 769 -1422
rect 833 -1456 867 -1422
rect 931 -1456 965 -1422
rect 1029 -1456 1063 -1422
rect 1127 -1456 1161 -1422
rect 1225 -1456 1259 -1422
rect 2204 160 2284 320
rect 2533 796 2567 830
rect 2631 796 2665 830
rect 2729 796 2763 830
rect 2827 796 2861 830
rect 2925 796 2959 830
rect 3023 796 3057 830
rect 3121 796 3155 830
rect 3219 796 3253 830
rect 3317 796 3351 830
rect 3415 796 3449 830
rect 3513 796 3547 830
rect 3611 796 3645 830
rect 3709 796 3743 830
rect 3807 796 3841 830
rect 3905 796 3939 830
rect 2484 370 2518 746
rect 2582 370 2616 746
rect 2680 370 2714 746
rect 2778 370 2812 746
rect 2876 370 2910 746
rect 2974 370 3008 746
rect 3072 370 3106 746
rect 3170 370 3204 746
rect 3268 370 3302 746
rect 3366 370 3400 746
rect 3464 370 3498 746
rect 3562 370 3596 746
rect 3660 370 3694 746
rect 3758 370 3792 746
rect 3856 370 3890 746
rect 3954 370 3988 746
rect 2533 286 2567 320
rect 2631 286 2665 320
rect 2729 286 2763 320
rect 2827 286 2861 320
rect 2925 286 2959 320
rect 3023 286 3057 320
rect 3121 286 3155 320
rect 3219 286 3253 320
rect 3317 286 3351 320
rect 3415 286 3449 320
rect 3513 286 3547 320
rect 3611 286 3645 320
rect 3709 286 3743 320
rect 3807 286 3841 320
rect 3905 286 3939 320
rect 2533 178 2567 212
rect 2631 178 2665 212
rect 2729 178 2763 212
rect 2827 178 2861 212
rect 2925 178 2959 212
rect 3023 178 3057 212
rect 3121 178 3155 212
rect 3219 178 3253 212
rect 3317 178 3351 212
rect 3415 178 3449 212
rect 3513 178 3547 212
rect 3611 178 3645 212
rect 3709 178 3743 212
rect 3807 178 3841 212
rect 3905 178 3939 212
rect 2484 -248 2518 128
rect 2582 -248 2616 128
rect 2680 -248 2714 128
rect 2778 -248 2812 128
rect 2876 -248 2910 128
rect 2974 -248 3008 128
rect 3072 -248 3106 128
rect 3170 -248 3204 128
rect 3268 -248 3302 128
rect 3366 -248 3400 128
rect 3464 -248 3498 128
rect 3562 -248 3596 128
rect 3660 -248 3694 128
rect 3758 -248 3792 128
rect 3856 -248 3890 128
rect 4054 130 4068 340
rect 4068 130 4102 340
rect 4102 130 4174 340
rect 3954 -248 3988 128
rect 2533 -332 2567 -298
rect 2631 -332 2665 -298
rect 2729 -332 2763 -298
rect 2827 -332 2861 -298
rect 2925 -332 2959 -298
rect 3023 -332 3057 -298
rect 3121 -332 3155 -298
rect 3219 -332 3253 -298
rect 3317 -332 3351 -298
rect 3415 -332 3449 -298
rect 3513 -332 3547 -298
rect 3611 -332 3645 -298
rect 3709 -332 3743 -298
rect 3807 -332 3841 -298
rect 3905 -332 3939 -298
rect 1662 -982 1696 -948
rect 1758 -982 1792 -948
rect 1854 -982 1888 -948
rect 1950 -982 1984 -948
rect 2046 -982 2080 -948
rect 2142 -982 2176 -948
rect 2238 -982 2272 -948
rect 2334 -982 2368 -948
rect 2430 -982 2464 -948
rect 2526 -982 2560 -948
rect 2622 -982 2656 -948
rect 2718 -982 2752 -948
rect 1614 -1408 1648 -1032
rect 1710 -1408 1744 -1032
rect 1806 -1408 1840 -1032
rect 1902 -1408 1936 -1032
rect 1998 -1408 2032 -1032
rect 2094 -1408 2128 -1032
rect 2190 -1408 2224 -1032
rect 2286 -1408 2320 -1032
rect 2382 -1408 2416 -1032
rect 2478 -1408 2512 -1032
rect 2574 -1408 2608 -1032
rect 2670 -1408 2704 -1032
rect 2766 -1408 2800 -1032
rect 1662 -1492 1696 -1458
rect 1758 -1492 1792 -1458
rect 1854 -1492 1888 -1458
rect 1950 -1492 1984 -1458
rect 2046 -1492 2080 -1458
rect 2142 -1492 2176 -1458
rect 2238 -1492 2272 -1458
rect 2334 -1492 2368 -1458
rect 2430 -1492 2464 -1458
rect 2526 -1492 2560 -1458
rect 2622 -1492 2656 -1458
rect 2718 -1492 2752 -1458
rect -1148 -1748 -1114 -1714
rect -956 -1748 -922 -1714
rect -764 -1748 -730 -1714
rect -572 -1748 -538 -1714
rect -380 -1748 -346 -1714
rect -188 -1748 -154 -1714
rect 4 -1748 38 -1714
rect 196 -1748 230 -1714
rect 388 -1748 422 -1714
rect 580 -1748 614 -1714
rect 772 -1748 806 -1714
rect 964 -1748 998 -1714
rect 1156 -1748 1190 -1714
rect -1196 -2174 -1162 -1798
rect -1100 -2174 -1066 -1798
rect -1004 -2174 -970 -1798
rect -908 -2174 -874 -1798
rect -812 -2174 -778 -1798
rect -716 -2174 -682 -1798
rect -620 -2174 -586 -1798
rect -524 -2174 -490 -1798
rect -428 -2174 -394 -1798
rect -332 -2174 -298 -1798
rect -236 -2174 -202 -1798
rect -140 -2174 -106 -1798
rect -44 -2174 -10 -1798
rect 52 -2174 86 -1798
rect 148 -2174 182 -1798
rect 244 -2174 278 -1798
rect 340 -2174 374 -1798
rect 436 -2174 470 -1798
rect 532 -2174 566 -1798
rect 628 -2174 662 -1798
rect 724 -2174 758 -1798
rect 820 -2174 854 -1798
rect 916 -2174 950 -1798
rect 1012 -2174 1046 -1798
rect 1108 -2174 1142 -1798
rect 1204 -2174 1238 -1798
rect -1052 -2258 -1018 -2224
rect -860 -2258 -826 -2224
rect -668 -2258 -634 -2224
rect -476 -2258 -442 -2224
rect -284 -2258 -250 -2224
rect -92 -2258 -58 -2224
rect 100 -2258 134 -2224
rect 292 -2258 326 -2224
rect 484 -2258 518 -2224
rect 676 -2258 710 -2224
rect 868 -2258 902 -2224
rect 1060 -2258 1094 -2224
rect 1344 -2250 1352 -2070
rect 1352 -2250 1474 -2070
rect -1052 -2366 -1018 -2332
rect -860 -2366 -826 -2332
rect -668 -2366 -634 -2332
rect -476 -2366 -442 -2332
rect -284 -2366 -250 -2332
rect -92 -2366 -58 -2332
rect 100 -2366 134 -2332
rect 292 -2366 326 -2332
rect 484 -2366 518 -2332
rect 676 -2366 710 -2332
rect 868 -2366 902 -2332
rect 1060 -2366 1094 -2332
rect -1196 -2792 -1162 -2416
rect -1100 -2792 -1066 -2416
rect -1004 -2792 -970 -2416
rect -908 -2792 -874 -2416
rect -812 -2792 -778 -2416
rect -716 -2792 -682 -2416
rect -620 -2792 -586 -2416
rect -524 -2792 -490 -2416
rect -428 -2792 -394 -2416
rect -332 -2792 -298 -2416
rect -236 -2792 -202 -2416
rect -140 -2792 -106 -2416
rect -44 -2792 -10 -2416
rect 52 -2792 86 -2416
rect 148 -2792 182 -2416
rect 244 -2792 278 -2416
rect 340 -2792 374 -2416
rect 436 -2792 470 -2416
rect 532 -2792 566 -2416
rect 628 -2792 662 -2416
rect 724 -2792 758 -2416
rect 820 -2792 854 -2416
rect 916 -2792 950 -2416
rect 1012 -2792 1046 -2416
rect 1108 -2792 1142 -2416
rect 1204 -2792 1238 -2416
rect -1148 -2876 -1114 -2842
rect -956 -2876 -922 -2842
rect -764 -2876 -730 -2842
rect -572 -2876 -538 -2842
rect -380 -2876 -346 -2842
rect -188 -2876 -154 -2842
rect 4 -2876 38 -2842
rect 196 -2876 230 -2842
rect 388 -2876 422 -2842
rect 580 -2876 614 -2842
rect 772 -2876 806 -2842
rect 964 -2876 998 -2842
rect 1156 -2876 1190 -2842
rect -1148 -2984 -1114 -2950
rect -956 -2984 -922 -2950
rect -764 -2984 -730 -2950
rect -572 -2984 -538 -2950
rect -380 -2984 -346 -2950
rect -188 -2984 -154 -2950
rect 4 -2984 38 -2950
rect 196 -2984 230 -2950
rect 388 -2984 422 -2950
rect 580 -2984 614 -2950
rect 772 -2984 806 -2950
rect 964 -2984 998 -2950
rect 1156 -2984 1190 -2950
rect -1196 -3410 -1162 -3034
rect -1100 -3410 -1066 -3034
rect -1004 -3410 -970 -3034
rect -908 -3410 -874 -3034
rect -812 -3410 -778 -3034
rect -716 -3410 -682 -3034
rect -620 -3410 -586 -3034
rect -524 -3410 -490 -3034
rect -428 -3410 -394 -3034
rect -332 -3410 -298 -3034
rect -236 -3410 -202 -3034
rect -140 -3410 -106 -3034
rect -44 -3410 -10 -3034
rect 52 -3410 86 -3034
rect 148 -3410 182 -3034
rect 244 -3410 278 -3034
rect 340 -3410 374 -3034
rect 436 -3410 470 -3034
rect 532 -3410 566 -3034
rect 628 -3410 662 -3034
rect 724 -3410 758 -3034
rect 820 -3410 854 -3034
rect 916 -3410 950 -3034
rect 1012 -3410 1046 -3034
rect 1108 -3410 1142 -3034
rect 1204 -3410 1238 -3034
rect -1052 -3494 -1018 -3460
rect -860 -3494 -826 -3460
rect -668 -3494 -634 -3460
rect -476 -3494 -442 -3460
rect -284 -3494 -250 -3460
rect -92 -3494 -58 -3460
rect 100 -3494 134 -3460
rect 292 -3494 326 -3460
rect 484 -3494 518 -3460
rect 676 -3494 710 -3460
rect 868 -3494 902 -3460
rect 1060 -3494 1094 -3460
rect -1052 -3602 -1018 -3568
rect -860 -3602 -826 -3568
rect -668 -3602 -634 -3568
rect -476 -3602 -442 -3568
rect -284 -3602 -250 -3568
rect -92 -3602 -58 -3568
rect 100 -3602 134 -3568
rect 292 -3602 326 -3568
rect 484 -3602 518 -3568
rect 676 -3602 710 -3568
rect 868 -3602 902 -3568
rect 1060 -3602 1094 -3568
rect -1196 -4028 -1162 -3652
rect -1100 -4028 -1066 -3652
rect -1004 -4028 -970 -3652
rect -908 -4028 -874 -3652
rect -812 -4028 -778 -3652
rect -716 -4028 -682 -3652
rect -620 -4028 -586 -3652
rect -524 -4028 -490 -3652
rect -428 -4028 -394 -3652
rect -332 -4028 -298 -3652
rect -236 -4028 -202 -3652
rect -140 -4028 -106 -3652
rect -44 -4028 -10 -3652
rect 52 -4028 86 -3652
rect 148 -4028 182 -3652
rect 244 -4028 278 -3652
rect 340 -4028 374 -3652
rect 436 -4028 470 -3652
rect 532 -4028 566 -3652
rect 628 -4028 662 -3652
rect 724 -4028 758 -3652
rect 820 -4028 854 -3652
rect 916 -4028 950 -3652
rect 1012 -4028 1046 -3652
rect 1108 -4028 1142 -3652
rect 1204 -4028 1238 -3652
rect -1148 -4112 -1114 -4078
rect -956 -4112 -922 -4078
rect -764 -4112 -730 -4078
rect -572 -4112 -538 -4078
rect -380 -4112 -346 -4078
rect -188 -4112 -154 -4078
rect 4 -4112 38 -4078
rect 196 -4112 230 -4078
rect 388 -4112 422 -4078
rect 580 -4112 614 -4078
rect 772 -4112 806 -4078
rect 964 -4112 998 -4078
rect 1156 -4112 1190 -4078
rect 1676 -1802 1844 -1768
rect 1934 -1802 2102 -1768
rect 2192 -1802 2360 -1768
rect 2450 -1802 2618 -1768
rect 2708 -1802 2876 -1768
rect 2966 -1802 3134 -1768
rect 1614 -2228 1648 -1852
rect 1872 -2228 1906 -1852
rect 2130 -2228 2164 -1852
rect 2388 -2228 2422 -1852
rect 2646 -2228 2680 -1852
rect 2904 -2228 2938 -1852
rect 3162 -2228 3196 -1852
rect 1676 -2312 1844 -2278
rect 1934 -2312 2102 -2278
rect 2192 -2312 2360 -2278
rect 2450 -2312 2618 -2278
rect 2708 -2312 2876 -2278
rect 2966 -2312 3134 -2278
rect -1127 -4478 -1093 -4444
rect -1029 -4478 -995 -4444
rect -931 -4478 -897 -4444
rect -833 -4478 -799 -4444
rect -735 -4478 -701 -4444
rect -637 -4478 -603 -4444
rect -539 -4478 -505 -4444
rect -441 -4478 -407 -4444
rect -343 -4478 -309 -4444
rect -245 -4478 -211 -4444
rect -147 -4478 -113 -4444
rect -49 -4478 -15 -4444
rect 49 -4478 83 -4444
rect 147 -4478 181 -4444
rect 245 -4478 279 -4444
rect -1176 -4913 -1142 -4537
rect -1078 -4913 -1044 -4537
rect -980 -4913 -946 -4537
rect -882 -4913 -848 -4537
rect -784 -4913 -750 -4537
rect -686 -4913 -652 -4537
rect -588 -4913 -554 -4537
rect -490 -4913 -456 -4537
rect -392 -4913 -358 -4537
rect -294 -4913 -260 -4537
rect -196 -4913 -162 -4537
rect -98 -4913 -64 -4537
rect 0 -4913 34 -4537
rect 98 -4913 132 -4537
rect 196 -4913 230 -4537
rect 294 -4913 328 -4537
rect -1127 -5006 -1093 -4972
rect -1029 -5006 -995 -4972
rect -931 -5006 -897 -4972
rect -833 -5006 -799 -4972
rect -735 -5006 -701 -4972
rect -637 -5006 -603 -4972
rect -539 -5006 -505 -4972
rect -441 -5006 -407 -4972
rect -343 -5006 -309 -4972
rect -245 -5006 -211 -4972
rect -147 -5006 -113 -4972
rect -49 -5006 -15 -4972
rect 49 -5006 83 -4972
rect 147 -5006 181 -4972
rect 245 -5006 279 -4972
rect -1127 -5114 -1093 -5080
rect -1029 -5114 -995 -5080
rect -931 -5114 -897 -5080
rect -833 -5114 -799 -5080
rect -735 -5114 -701 -5080
rect -637 -5114 -603 -5080
rect -539 -5114 -505 -5080
rect -441 -5114 -407 -5080
rect -343 -5114 -309 -5080
rect -245 -5114 -211 -5080
rect -147 -5114 -113 -5080
rect -49 -5114 -15 -5080
rect 49 -5114 83 -5080
rect 147 -5114 181 -5080
rect 245 -5114 279 -5080
rect -1176 -5549 -1142 -5173
rect -1078 -5549 -1044 -5173
rect -980 -5549 -946 -5173
rect -882 -5549 -848 -5173
rect -784 -5549 -750 -5173
rect -686 -5549 -652 -5173
rect -588 -5549 -554 -5173
rect -490 -5549 -456 -5173
rect -392 -5549 -358 -5173
rect -294 -5549 -260 -5173
rect -196 -5549 -162 -5173
rect -98 -5549 -64 -5173
rect 0 -5549 34 -5173
rect 98 -5549 132 -5173
rect 196 -5549 230 -5173
rect 294 -5549 328 -5173
rect -1127 -5642 -1093 -5608
rect -1029 -5642 -995 -5608
rect -931 -5642 -897 -5608
rect -833 -5642 -799 -5608
rect -735 -5642 -701 -5608
rect -637 -5642 -603 -5608
rect -539 -5642 -505 -5608
rect -441 -5642 -407 -5608
rect -343 -5642 -309 -5608
rect -245 -5642 -211 -5608
rect -147 -5642 -113 -5608
rect -49 -5642 -15 -5608
rect 49 -5642 83 -5608
rect 147 -5642 181 -5608
rect 245 -5642 279 -5608
rect 671 -4478 705 -4444
rect 769 -4478 803 -4444
rect 867 -4478 901 -4444
rect 965 -4478 999 -4444
rect 1063 -4478 1097 -4444
rect 1161 -4478 1195 -4444
rect 1259 -4478 1293 -4444
rect 1357 -4478 1391 -4444
rect 1455 -4478 1489 -4444
rect 1553 -4478 1587 -4444
rect 1651 -4478 1685 -4444
rect 1749 -4478 1783 -4444
rect 1847 -4478 1881 -4444
rect 1945 -4478 1979 -4444
rect 2043 -4478 2077 -4444
rect 622 -4913 656 -4537
rect 720 -4913 754 -4537
rect 818 -4913 852 -4537
rect 916 -4913 950 -4537
rect 1014 -4913 1048 -4537
rect 1112 -4913 1146 -4537
rect 1210 -4913 1244 -4537
rect 1308 -4913 1342 -4537
rect 1406 -4913 1440 -4537
rect 1504 -4913 1538 -4537
rect 1602 -4913 1636 -4537
rect 1700 -4913 1734 -4537
rect 1798 -4913 1832 -4537
rect 1896 -4913 1930 -4537
rect 1994 -4913 2028 -4537
rect 2092 -4913 2126 -4537
rect 671 -5006 705 -4972
rect 769 -5006 803 -4972
rect 867 -5006 901 -4972
rect 965 -5006 999 -4972
rect 1063 -5006 1097 -4972
rect 1161 -5006 1195 -4972
rect 1259 -5006 1293 -4972
rect 1357 -5006 1391 -4972
rect 1455 -5006 1489 -4972
rect 1553 -5006 1587 -4972
rect 1651 -5006 1685 -4972
rect 1749 -5006 1783 -4972
rect 1847 -5006 1881 -4972
rect 1945 -5006 1979 -4972
rect 2043 -5006 2077 -4972
rect 671 -5114 705 -5080
rect 769 -5114 803 -5080
rect 867 -5114 901 -5080
rect 965 -5114 999 -5080
rect 1063 -5114 1097 -5080
rect 1161 -5114 1195 -5080
rect 1259 -5114 1293 -5080
rect 1357 -5114 1391 -5080
rect 1455 -5114 1489 -5080
rect 1553 -5114 1587 -5080
rect 1651 -5114 1685 -5080
rect 1749 -5114 1783 -5080
rect 1847 -5114 1881 -5080
rect 1945 -5114 1979 -5080
rect 2043 -5114 2077 -5080
rect 622 -5549 656 -5173
rect 720 -5549 754 -5173
rect 818 -5549 852 -5173
rect 916 -5549 950 -5173
rect 1014 -5549 1048 -5173
rect 1112 -5549 1146 -5173
rect 1210 -5549 1244 -5173
rect 1308 -5549 1342 -5173
rect 1406 -5549 1440 -5173
rect 1504 -5549 1538 -5173
rect 1602 -5549 1636 -5173
rect 1700 -5549 1734 -5173
rect 1798 -5549 1832 -5173
rect 1896 -5549 1930 -5173
rect 1994 -5549 2028 -5173
rect 2092 -5549 2126 -5173
rect 2214 -5560 2240 -5000
rect 2240 -5090 2344 -5000
rect 2240 -5560 2310 -5090
rect 2310 -5560 2344 -5090
rect 2486 -5130 2554 -5096
rect 2644 -5130 2712 -5096
rect 2802 -5130 2870 -5096
rect 2960 -5130 3028 -5096
rect 3118 -5130 3186 -5096
rect 3276 -5130 3344 -5096
rect 3434 -5130 3502 -5096
rect 3592 -5130 3660 -5096
rect 3750 -5130 3818 -5096
rect 3908 -5130 3976 -5096
rect 671 -5642 705 -5608
rect 769 -5642 803 -5608
rect 867 -5642 901 -5608
rect 965 -5642 999 -5608
rect 1063 -5642 1097 -5608
rect 1161 -5642 1195 -5608
rect 1259 -5642 1293 -5608
rect 1357 -5642 1391 -5608
rect 1455 -5642 1489 -5608
rect 1553 -5642 1587 -5608
rect 1651 -5642 1685 -5608
rect 1749 -5642 1783 -5608
rect 1847 -5642 1881 -5608
rect 1945 -5642 1979 -5608
rect 2043 -5642 2077 -5608
rect 2424 -5565 2458 -5189
rect 2582 -5565 2616 -5189
rect 2740 -5565 2774 -5189
rect 2898 -5565 2932 -5189
rect 3056 -5565 3090 -5189
rect 3214 -5565 3248 -5189
rect 3372 -5565 3406 -5189
rect 3530 -5565 3564 -5189
rect 3688 -5565 3722 -5189
rect 3846 -5565 3880 -5189
rect 4004 -5565 4038 -5189
rect 2486 -5658 2554 -5624
rect 2644 -5658 2712 -5624
rect 2802 -5658 2870 -5624
rect 2960 -5658 3028 -5624
rect 3118 -5658 3186 -5624
rect 3276 -5658 3344 -5624
rect 3434 -5658 3502 -5624
rect 3592 -5658 3660 -5624
rect 3750 -5658 3818 -5624
rect 3908 -5658 3976 -5624
rect -1127 -5954 -1093 -5920
rect -1030 -5954 -996 -5920
rect -931 -5954 -897 -5920
rect -834 -5954 -800 -5920
rect -735 -5954 -701 -5920
rect -638 -5954 -604 -5920
rect -539 -5954 -505 -5920
rect -442 -5954 -408 -5920
rect -343 -5954 -309 -5920
rect -246 -5954 -212 -5920
rect -147 -5954 -113 -5920
rect -50 -5954 -16 -5920
rect 49 -5954 83 -5920
rect 146 -5954 180 -5920
rect 245 -5954 279 -5920
rect 342 -5954 376 -5920
rect 441 -5954 475 -5920
rect 538 -5954 572 -5920
rect 637 -5954 671 -5920
rect 734 -5954 768 -5920
rect 833 -5954 867 -5920
rect 930 -5954 964 -5920
rect 1029 -5954 1063 -5920
rect 1126 -5954 1160 -5920
rect 1225 -5954 1259 -5920
rect -1176 -6380 -1142 -6004
rect -1078 -6380 -1044 -6004
rect -980 -6380 -946 -6004
rect -882 -6380 -848 -6004
rect -784 -6380 -750 -6004
rect -686 -6380 -652 -6004
rect -588 -6380 -554 -6004
rect -490 -6380 -456 -6004
rect -392 -6380 -358 -6004
rect -294 -6380 -260 -6004
rect -196 -6380 -162 -6004
rect -98 -6380 -64 -6004
rect 0 -6380 34 -6004
rect 98 -6380 132 -6004
rect 196 -6380 230 -6004
rect 294 -6380 328 -6004
rect 392 -6380 426 -6004
rect 490 -6380 524 -6004
rect 588 -6380 622 -6004
rect 686 -6380 720 -6004
rect 784 -6380 818 -6004
rect 882 -6380 916 -6004
rect 980 -6380 1014 -6004
rect 1078 -6380 1112 -6004
rect 1176 -6380 1210 -6004
rect 1274 -6380 1308 -6004
rect -1128 -6464 -1094 -6430
rect -1029 -6464 -995 -6430
rect -932 -6464 -898 -6430
rect -833 -6464 -799 -6430
rect -736 -6464 -702 -6430
rect -637 -6464 -603 -6430
rect -540 -6464 -506 -6430
rect -441 -6464 -407 -6430
rect -344 -6464 -310 -6430
rect -245 -6464 -211 -6430
rect -148 -6464 -114 -6430
rect -49 -6464 -15 -6430
rect 48 -6464 82 -6430
rect 147 -6464 181 -6430
rect 244 -6464 278 -6430
rect 343 -6464 377 -6430
rect 440 -6464 474 -6430
rect 539 -6464 573 -6430
rect 636 -6464 670 -6430
rect 735 -6464 769 -6430
rect 832 -6464 866 -6430
rect 931 -6464 965 -6430
rect 1028 -6464 1062 -6430
rect 1127 -6464 1161 -6430
rect 1224 -6464 1258 -6430
rect -1127 -6572 -1093 -6538
rect -1029 -6572 -995 -6538
rect -931 -6572 -897 -6538
rect -833 -6572 -799 -6538
rect -735 -6572 -701 -6538
rect -637 -6572 -603 -6538
rect -539 -6572 -505 -6538
rect -441 -6572 -407 -6538
rect -343 -6572 -309 -6538
rect -245 -6572 -211 -6538
rect -147 -6572 -113 -6538
rect -49 -6572 -15 -6538
rect 49 -6572 83 -6538
rect 147 -6572 181 -6538
rect 245 -6572 279 -6538
rect 343 -6572 377 -6538
rect 441 -6572 475 -6538
rect 539 -6572 573 -6538
rect 637 -6572 671 -6538
rect 735 -6572 769 -6538
rect 833 -6572 867 -6538
rect 931 -6572 965 -6538
rect 1029 -6572 1063 -6538
rect 1127 -6572 1161 -6538
rect 1225 -6572 1259 -6538
rect -1176 -6998 -1142 -6622
rect -1078 -6998 -1044 -6622
rect -980 -6998 -946 -6622
rect -882 -6998 -848 -6622
rect -784 -6998 -750 -6622
rect -686 -6998 -652 -6622
rect -588 -6998 -554 -6622
rect -490 -6998 -456 -6622
rect -392 -6998 -358 -6622
rect -294 -6998 -260 -6622
rect -196 -6998 -162 -6622
rect -98 -6998 -64 -6622
rect 0 -6998 34 -6622
rect 98 -6998 132 -6622
rect 196 -6998 230 -6622
rect 294 -6998 328 -6622
rect 392 -6998 426 -6622
rect 490 -6998 524 -6622
rect 588 -6998 622 -6622
rect 686 -6998 720 -6622
rect 784 -6998 818 -6622
rect 882 -6998 916 -6622
rect 980 -6998 1014 -6622
rect 1078 -6998 1112 -6622
rect 1176 -6998 1210 -6622
rect 1274 -6998 1308 -6622
rect -1127 -7082 -1093 -7048
rect -1029 -7082 -995 -7048
rect -931 -7082 -897 -7048
rect -833 -7082 -799 -7048
rect -735 -7082 -701 -7048
rect -637 -7082 -603 -7048
rect -539 -7082 -505 -7048
rect -441 -7082 -407 -7048
rect -343 -7082 -309 -7048
rect -245 -7082 -211 -7048
rect -147 -7082 -113 -7048
rect -49 -7082 -15 -7048
rect 49 -7082 83 -7048
rect 147 -7082 181 -7048
rect 245 -7082 279 -7048
rect 343 -7082 377 -7048
rect 441 -7082 475 -7048
rect 539 -7082 573 -7048
rect 637 -7082 671 -7048
rect 735 -7082 769 -7048
rect 833 -7082 867 -7048
rect 931 -7082 965 -7048
rect 1029 -7082 1063 -7048
rect 1127 -7082 1161 -7048
rect 1225 -7082 1259 -7048
rect -1127 -7398 -1093 -7364
rect -1030 -7398 -996 -7364
rect -931 -7398 -897 -7364
rect -834 -7398 -800 -7364
rect -735 -7398 -701 -7364
rect -638 -7398 -604 -7364
rect -539 -7398 -505 -7364
rect -442 -7398 -408 -7364
rect -343 -7398 -309 -7364
rect -246 -7398 -212 -7364
rect -147 -7398 -113 -7364
rect -50 -7398 -16 -7364
rect 49 -7398 83 -7364
rect 146 -7398 180 -7364
rect 245 -7398 279 -7364
rect 342 -7398 376 -7364
rect 441 -7398 475 -7364
rect 538 -7398 572 -7364
rect 637 -7398 671 -7364
rect 734 -7398 768 -7364
rect 833 -7398 867 -7364
rect 930 -7398 964 -7364
rect 1029 -7398 1063 -7364
rect 1126 -7398 1160 -7364
rect 1225 -7398 1259 -7364
rect -1176 -7824 -1142 -7448
rect -1078 -7824 -1044 -7448
rect -980 -7824 -946 -7448
rect -882 -7824 -848 -7448
rect -784 -7824 -750 -7448
rect -686 -7824 -652 -7448
rect -588 -7824 -554 -7448
rect -490 -7824 -456 -7448
rect -392 -7824 -358 -7448
rect -294 -7824 -260 -7448
rect -196 -7824 -162 -7448
rect -98 -7824 -64 -7448
rect 0 -7824 34 -7448
rect 98 -7824 132 -7448
rect 196 -7824 230 -7448
rect 294 -7824 328 -7448
rect 392 -7824 426 -7448
rect 490 -7824 524 -7448
rect 588 -7824 622 -7448
rect 686 -7824 720 -7448
rect 784 -7824 818 -7448
rect 882 -7824 916 -7448
rect 980 -7824 1014 -7448
rect 1078 -7824 1112 -7448
rect 1176 -7824 1210 -7448
rect 1274 -7824 1308 -7448
rect -1128 -7908 -1094 -7874
rect -1029 -7908 -995 -7874
rect -932 -7908 -898 -7874
rect -833 -7908 -799 -7874
rect -736 -7908 -702 -7874
rect -637 -7908 -603 -7874
rect -540 -7908 -506 -7874
rect -441 -7908 -407 -7874
rect -344 -7908 -310 -7874
rect -245 -7908 -211 -7874
rect -148 -7908 -114 -7874
rect -49 -7908 -15 -7874
rect 48 -7908 82 -7874
rect 147 -7908 181 -7874
rect 244 -7908 278 -7874
rect 343 -7908 377 -7874
rect 440 -7908 474 -7874
rect 539 -7908 573 -7874
rect 636 -7908 670 -7874
rect 735 -7908 769 -7874
rect 832 -7908 866 -7874
rect 931 -7908 965 -7874
rect 1028 -7908 1062 -7874
rect 1127 -7908 1161 -7874
rect 1224 -7908 1258 -7874
rect -1127 -8016 -1093 -7982
rect -1029 -8016 -995 -7982
rect -931 -8016 -897 -7982
rect -833 -8016 -799 -7982
rect -735 -8016 -701 -7982
rect -637 -8016 -603 -7982
rect -539 -8016 -505 -7982
rect -441 -8016 -407 -7982
rect -343 -8016 -309 -7982
rect -245 -8016 -211 -7982
rect -147 -8016 -113 -7982
rect -49 -8016 -15 -7982
rect 49 -8016 83 -7982
rect 147 -8016 181 -7982
rect 245 -8016 279 -7982
rect 343 -8016 377 -7982
rect 441 -8016 475 -7982
rect 539 -8016 573 -7982
rect 637 -8016 671 -7982
rect 735 -8016 769 -7982
rect 833 -8016 867 -7982
rect 931 -8016 965 -7982
rect 1029 -8016 1063 -7982
rect 1127 -8016 1161 -7982
rect 1225 -8016 1259 -7982
rect -1176 -8442 -1142 -8066
rect -1078 -8442 -1044 -8066
rect -980 -8442 -946 -8066
rect -882 -8442 -848 -8066
rect -784 -8442 -750 -8066
rect -686 -8442 -652 -8066
rect -588 -8442 -554 -8066
rect -490 -8442 -456 -8066
rect -392 -8442 -358 -8066
rect -294 -8442 -260 -8066
rect -196 -8442 -162 -8066
rect -98 -8442 -64 -8066
rect 0 -8442 34 -8066
rect 98 -8442 132 -8066
rect 196 -8442 230 -8066
rect 294 -8442 328 -8066
rect 392 -8442 426 -8066
rect 490 -8442 524 -8066
rect 588 -8442 622 -8066
rect 686 -8442 720 -8066
rect 784 -8442 818 -8066
rect 882 -8442 916 -8066
rect 980 -8442 1014 -8066
rect 1078 -8442 1112 -8066
rect 1176 -8442 1210 -8066
rect 1274 -8442 1308 -8066
rect -1127 -8526 -1093 -8492
rect -1029 -8526 -995 -8492
rect -931 -8526 -897 -8492
rect -833 -8526 -799 -8492
rect -735 -8526 -701 -8492
rect -637 -8526 -603 -8492
rect -539 -8526 -505 -8492
rect -441 -8526 -407 -8492
rect -343 -8526 -309 -8492
rect -245 -8526 -211 -8492
rect -147 -8526 -113 -8492
rect -49 -8526 -15 -8492
rect 49 -8526 83 -8492
rect 147 -8526 181 -8492
rect 245 -8526 279 -8492
rect 343 -8526 377 -8492
rect 441 -8526 475 -8492
rect 539 -8526 573 -8492
rect 637 -8526 671 -8492
rect 735 -8526 769 -8492
rect 833 -8526 867 -8492
rect 931 -8526 965 -8492
rect 1029 -8526 1063 -8492
rect 1127 -8526 1161 -8492
rect 1225 -8526 1259 -8492
rect 2204 -6910 2284 -6750
rect 2533 -6274 2567 -6240
rect 2631 -6274 2665 -6240
rect 2729 -6274 2763 -6240
rect 2827 -6274 2861 -6240
rect 2925 -6274 2959 -6240
rect 3023 -6274 3057 -6240
rect 3121 -6274 3155 -6240
rect 3219 -6274 3253 -6240
rect 3317 -6274 3351 -6240
rect 3415 -6274 3449 -6240
rect 3513 -6274 3547 -6240
rect 3611 -6274 3645 -6240
rect 3709 -6274 3743 -6240
rect 3807 -6274 3841 -6240
rect 3905 -6274 3939 -6240
rect 2484 -6700 2518 -6324
rect 2582 -6700 2616 -6324
rect 2680 -6700 2714 -6324
rect 2778 -6700 2812 -6324
rect 2876 -6700 2910 -6324
rect 2974 -6700 3008 -6324
rect 3072 -6700 3106 -6324
rect 3170 -6700 3204 -6324
rect 3268 -6700 3302 -6324
rect 3366 -6700 3400 -6324
rect 3464 -6700 3498 -6324
rect 3562 -6700 3596 -6324
rect 3660 -6700 3694 -6324
rect 3758 -6700 3792 -6324
rect 3856 -6700 3890 -6324
rect 3954 -6700 3988 -6324
rect 2533 -6784 2567 -6750
rect 2631 -6784 2665 -6750
rect 2729 -6784 2763 -6750
rect 2827 -6784 2861 -6750
rect 2925 -6784 2959 -6750
rect 3023 -6784 3057 -6750
rect 3121 -6784 3155 -6750
rect 3219 -6784 3253 -6750
rect 3317 -6784 3351 -6750
rect 3415 -6784 3449 -6750
rect 3513 -6784 3547 -6750
rect 3611 -6784 3645 -6750
rect 3709 -6784 3743 -6750
rect 3807 -6784 3841 -6750
rect 3905 -6784 3939 -6750
rect 2533 -6892 2567 -6858
rect 2631 -6892 2665 -6858
rect 2729 -6892 2763 -6858
rect 2827 -6892 2861 -6858
rect 2925 -6892 2959 -6858
rect 3023 -6892 3057 -6858
rect 3121 -6892 3155 -6858
rect 3219 -6892 3253 -6858
rect 3317 -6892 3351 -6858
rect 3415 -6892 3449 -6858
rect 3513 -6892 3547 -6858
rect 3611 -6892 3645 -6858
rect 3709 -6892 3743 -6858
rect 3807 -6892 3841 -6858
rect 3905 -6892 3939 -6858
rect 2484 -7318 2518 -6942
rect 2582 -7318 2616 -6942
rect 2680 -7318 2714 -6942
rect 2778 -7318 2812 -6942
rect 2876 -7318 2910 -6942
rect 2974 -7318 3008 -6942
rect 3072 -7318 3106 -6942
rect 3170 -7318 3204 -6942
rect 3268 -7318 3302 -6942
rect 3366 -7318 3400 -6942
rect 3464 -7318 3498 -6942
rect 3562 -7318 3596 -6942
rect 3660 -7318 3694 -6942
rect 3758 -7318 3792 -6942
rect 3856 -7318 3890 -6942
rect 4054 -6940 4068 -6730
rect 4068 -6940 4102 -6730
rect 4102 -6940 4174 -6730
rect 3954 -7318 3988 -6942
rect 2533 -7402 2567 -7368
rect 2631 -7402 2665 -7368
rect 2729 -7402 2763 -7368
rect 2827 -7402 2861 -7368
rect 2925 -7402 2959 -7368
rect 3023 -7402 3057 -7368
rect 3121 -7402 3155 -7368
rect 3219 -7402 3253 -7368
rect 3317 -7402 3351 -7368
rect 3415 -7402 3449 -7368
rect 3513 -7402 3547 -7368
rect 3611 -7402 3645 -7368
rect 3709 -7402 3743 -7368
rect 3807 -7402 3841 -7368
rect 3905 -7402 3939 -7368
rect 1662 -8052 1696 -8018
rect 1758 -8052 1792 -8018
rect 1854 -8052 1888 -8018
rect 1950 -8052 1984 -8018
rect 2046 -8052 2080 -8018
rect 2142 -8052 2176 -8018
rect 2238 -8052 2272 -8018
rect 2334 -8052 2368 -8018
rect 2430 -8052 2464 -8018
rect 2526 -8052 2560 -8018
rect 2622 -8052 2656 -8018
rect 2718 -8052 2752 -8018
rect 1614 -8478 1648 -8102
rect 1710 -8478 1744 -8102
rect 1806 -8478 1840 -8102
rect 1902 -8478 1936 -8102
rect 1998 -8478 2032 -8102
rect 2094 -8478 2128 -8102
rect 2190 -8478 2224 -8102
rect 2286 -8478 2320 -8102
rect 2382 -8478 2416 -8102
rect 2478 -8478 2512 -8102
rect 2574 -8478 2608 -8102
rect 2670 -8478 2704 -8102
rect 2766 -8478 2800 -8102
rect 1662 -8562 1696 -8528
rect 1758 -8562 1792 -8528
rect 1854 -8562 1888 -8528
rect 1950 -8562 1984 -8528
rect 2046 -8562 2080 -8528
rect 2142 -8562 2176 -8528
rect 2238 -8562 2272 -8528
rect 2334 -8562 2368 -8528
rect 2430 -8562 2464 -8528
rect 2526 -8562 2560 -8528
rect 2622 -8562 2656 -8528
rect 2718 -8562 2752 -8528
rect 3558 -8052 3592 -8018
rect 3654 -8052 3688 -8018
rect 3750 -8052 3784 -8018
rect 3846 -8052 3880 -8018
rect 3942 -8052 3976 -8018
rect 4038 -8052 4072 -8018
rect 4134 -8052 4168 -8018
rect 4230 -8052 4264 -8018
rect 4326 -8052 4360 -8018
rect 4422 -8052 4456 -8018
rect 4518 -8052 4552 -8018
rect 4614 -8052 4648 -8018
rect 3510 -8478 3544 -8102
rect 3606 -8478 3640 -8102
rect 3702 -8478 3736 -8102
rect 3798 -8478 3832 -8102
rect 3894 -8478 3928 -8102
rect 3990 -8478 4024 -8102
rect 4086 -8478 4120 -8102
rect 4182 -8478 4216 -8102
rect 4278 -8478 4312 -8102
rect 4374 -8478 4408 -8102
rect 4470 -8478 4504 -8102
rect 4566 -8478 4600 -8102
rect 4662 -8478 4696 -8102
rect 3558 -8562 3592 -8528
rect 3654 -8562 3688 -8528
rect 3750 -8562 3784 -8528
rect 3846 -8562 3880 -8528
rect 3942 -8562 3976 -8528
rect 4038 -8562 4072 -8528
rect 4134 -8562 4168 -8528
rect 4230 -8562 4264 -8528
rect 4326 -8562 4360 -8528
rect 4422 -8562 4456 -8528
rect 4518 -8562 4552 -8528
rect 4614 -8562 4648 -8528
rect -1148 -8818 -1114 -8784
rect -956 -8818 -922 -8784
rect -764 -8818 -730 -8784
rect -572 -8818 -538 -8784
rect -380 -8818 -346 -8784
rect -188 -8818 -154 -8784
rect 4 -8818 38 -8784
rect 196 -8818 230 -8784
rect 388 -8818 422 -8784
rect 580 -8818 614 -8784
rect 772 -8818 806 -8784
rect 964 -8818 998 -8784
rect 1156 -8818 1190 -8784
rect -1196 -9244 -1162 -8868
rect -1100 -9244 -1066 -8868
rect -1004 -9244 -970 -8868
rect -908 -9244 -874 -8868
rect -812 -9244 -778 -8868
rect -716 -9244 -682 -8868
rect -620 -9244 -586 -8868
rect -524 -9244 -490 -8868
rect -428 -9244 -394 -8868
rect -332 -9244 -298 -8868
rect -236 -9244 -202 -8868
rect -140 -9244 -106 -8868
rect -44 -9244 -10 -8868
rect 52 -9244 86 -8868
rect 148 -9244 182 -8868
rect 244 -9244 278 -8868
rect 340 -9244 374 -8868
rect 436 -9244 470 -8868
rect 532 -9244 566 -8868
rect 628 -9244 662 -8868
rect 724 -9244 758 -8868
rect 820 -9244 854 -8868
rect 916 -9244 950 -8868
rect 1012 -9244 1046 -8868
rect 1108 -9244 1142 -8868
rect 1204 -9244 1238 -8868
rect -1052 -9328 -1018 -9294
rect -860 -9328 -826 -9294
rect -668 -9328 -634 -9294
rect -476 -9328 -442 -9294
rect -284 -9328 -250 -9294
rect -92 -9328 -58 -9294
rect 100 -9328 134 -9294
rect 292 -9328 326 -9294
rect 484 -9328 518 -9294
rect 676 -9328 710 -9294
rect 868 -9328 902 -9294
rect 1060 -9328 1094 -9294
rect 1344 -9320 1352 -9140
rect 1352 -9320 1474 -9140
rect -1052 -9436 -1018 -9402
rect -860 -9436 -826 -9402
rect -668 -9436 -634 -9402
rect -476 -9436 -442 -9402
rect -284 -9436 -250 -9402
rect -92 -9436 -58 -9402
rect 100 -9436 134 -9402
rect 292 -9436 326 -9402
rect 484 -9436 518 -9402
rect 676 -9436 710 -9402
rect 868 -9436 902 -9402
rect 1060 -9436 1094 -9402
rect -1196 -9862 -1162 -9486
rect -1100 -9862 -1066 -9486
rect -1004 -9862 -970 -9486
rect -908 -9862 -874 -9486
rect -812 -9862 -778 -9486
rect -716 -9862 -682 -9486
rect -620 -9862 -586 -9486
rect -524 -9862 -490 -9486
rect -428 -9862 -394 -9486
rect -332 -9862 -298 -9486
rect -236 -9862 -202 -9486
rect -140 -9862 -106 -9486
rect -44 -9862 -10 -9486
rect 52 -9862 86 -9486
rect 148 -9862 182 -9486
rect 244 -9862 278 -9486
rect 340 -9862 374 -9486
rect 436 -9862 470 -9486
rect 532 -9862 566 -9486
rect 628 -9862 662 -9486
rect 724 -9862 758 -9486
rect 820 -9862 854 -9486
rect 916 -9862 950 -9486
rect 1012 -9862 1046 -9486
rect 1108 -9862 1142 -9486
rect 1204 -9862 1238 -9486
rect -1148 -9946 -1114 -9912
rect -956 -9946 -922 -9912
rect -764 -9946 -730 -9912
rect -572 -9946 -538 -9912
rect -380 -9946 -346 -9912
rect -188 -9946 -154 -9912
rect 4 -9946 38 -9912
rect 196 -9946 230 -9912
rect 388 -9946 422 -9912
rect 580 -9946 614 -9912
rect 772 -9946 806 -9912
rect 964 -9946 998 -9912
rect 1156 -9946 1190 -9912
rect -1148 -10054 -1114 -10020
rect -956 -10054 -922 -10020
rect -764 -10054 -730 -10020
rect -572 -10054 -538 -10020
rect -380 -10054 -346 -10020
rect -188 -10054 -154 -10020
rect 4 -10054 38 -10020
rect 196 -10054 230 -10020
rect 388 -10054 422 -10020
rect 580 -10054 614 -10020
rect 772 -10054 806 -10020
rect 964 -10054 998 -10020
rect 1156 -10054 1190 -10020
rect -1196 -10480 -1162 -10104
rect -1100 -10480 -1066 -10104
rect -1004 -10480 -970 -10104
rect -908 -10480 -874 -10104
rect -812 -10480 -778 -10104
rect -716 -10480 -682 -10104
rect -620 -10480 -586 -10104
rect -524 -10480 -490 -10104
rect -428 -10480 -394 -10104
rect -332 -10480 -298 -10104
rect -236 -10480 -202 -10104
rect -140 -10480 -106 -10104
rect -44 -10480 -10 -10104
rect 52 -10480 86 -10104
rect 148 -10480 182 -10104
rect 244 -10480 278 -10104
rect 340 -10480 374 -10104
rect 436 -10480 470 -10104
rect 532 -10480 566 -10104
rect 628 -10480 662 -10104
rect 724 -10480 758 -10104
rect 820 -10480 854 -10104
rect 916 -10480 950 -10104
rect 1012 -10480 1046 -10104
rect 1108 -10480 1142 -10104
rect 1204 -10480 1238 -10104
rect -1052 -10564 -1018 -10530
rect -860 -10564 -826 -10530
rect -668 -10564 -634 -10530
rect -476 -10564 -442 -10530
rect -284 -10564 -250 -10530
rect -92 -10564 -58 -10530
rect 100 -10564 134 -10530
rect 292 -10564 326 -10530
rect 484 -10564 518 -10530
rect 676 -10564 710 -10530
rect 868 -10564 902 -10530
rect 1060 -10564 1094 -10530
rect -1052 -10672 -1018 -10638
rect -860 -10672 -826 -10638
rect -668 -10672 -634 -10638
rect -476 -10672 -442 -10638
rect -284 -10672 -250 -10638
rect -92 -10672 -58 -10638
rect 100 -10672 134 -10638
rect 292 -10672 326 -10638
rect 484 -10672 518 -10638
rect 676 -10672 710 -10638
rect 868 -10672 902 -10638
rect 1060 -10672 1094 -10638
rect -1196 -11098 -1162 -10722
rect -1100 -11098 -1066 -10722
rect -1004 -11098 -970 -10722
rect -908 -11098 -874 -10722
rect -812 -11098 -778 -10722
rect -716 -11098 -682 -10722
rect -620 -11098 -586 -10722
rect -524 -11098 -490 -10722
rect -428 -11098 -394 -10722
rect -332 -11098 -298 -10722
rect -236 -11098 -202 -10722
rect -140 -11098 -106 -10722
rect -44 -11098 -10 -10722
rect 52 -11098 86 -10722
rect 148 -11098 182 -10722
rect 244 -11098 278 -10722
rect 340 -11098 374 -10722
rect 436 -11098 470 -10722
rect 532 -11098 566 -10722
rect 628 -11098 662 -10722
rect 724 -11098 758 -10722
rect 820 -11098 854 -10722
rect 916 -11098 950 -10722
rect 1012 -11098 1046 -10722
rect 1108 -11098 1142 -10722
rect 1204 -11098 1238 -10722
rect -1148 -11182 -1114 -11148
rect -956 -11182 -922 -11148
rect -764 -11182 -730 -11148
rect -572 -11182 -538 -11148
rect -380 -11182 -346 -11148
rect -188 -11182 -154 -11148
rect 4 -11182 38 -11148
rect 196 -11182 230 -11148
rect 388 -11182 422 -11148
rect 580 -11182 614 -11148
rect 772 -11182 806 -11148
rect 964 -11182 998 -11148
rect 1156 -11182 1190 -11148
rect 1676 -8872 1844 -8838
rect 1934 -8872 2102 -8838
rect 2192 -8872 2360 -8838
rect 2450 -8872 2618 -8838
rect 2708 -8872 2876 -8838
rect 2966 -8872 3134 -8838
rect 1614 -9298 1648 -8922
rect 1872 -9298 1906 -8922
rect 2130 -9298 2164 -8922
rect 2388 -9298 2422 -8922
rect 2646 -9298 2680 -8922
rect 2904 -9298 2938 -8922
rect 3162 -9298 3196 -8922
rect 1676 -9382 1844 -9348
rect 1934 -9382 2102 -9348
rect 2192 -9382 2360 -9348
rect 2450 -9382 2618 -9348
rect 2708 -9382 2876 -9348
rect 2966 -9382 3134 -9348
rect 3572 -8872 3740 -8838
rect 3830 -8872 3998 -8838
rect 4088 -8872 4256 -8838
rect 4346 -8872 4514 -8838
rect 4604 -8872 4772 -8838
rect 4862 -8872 5030 -8838
rect 3510 -9298 3544 -8922
rect 3768 -9298 3802 -8922
rect 4026 -9298 4060 -8922
rect 4284 -9298 4318 -8922
rect 4542 -9298 4576 -8922
rect 4800 -9298 4834 -8922
rect 5058 -9298 5092 -8922
rect 3572 -9382 3740 -9348
rect 3830 -9382 3998 -9348
rect 4088 -9382 4256 -9348
rect 4346 -9382 4514 -9348
rect 4604 -9382 4772 -9348
rect 4862 -9382 5030 -9348
rect 5604 -8872 5638 -8838
rect 5796 -8872 5830 -8838
rect 5460 -9298 5494 -8922
rect 5556 -9298 5590 -8922
rect 5652 -9298 5686 -8922
rect 5748 -9298 5782 -8922
rect 5844 -9298 5878 -8922
rect 5940 -9298 5974 -8922
rect 5508 -9382 5542 -9348
rect 5700 -9382 5734 -9348
rect 5892 -9382 5926 -9348
rect 1709 -9884 2077 -9850
rect 2629 -9884 2997 -9850
rect 3549 -9884 3917 -9850
rect 4469 -9884 4837 -9850
rect 5389 -9884 5757 -9850
rect 1608 -10898 1642 -9946
rect 2144 -10898 2178 -9946
rect 2528 -10898 2562 -9946
rect 3064 -10898 3098 -9946
rect 3448 -10898 3482 -9946
rect 3984 -10898 4018 -9946
rect 4368 -10898 4402 -9946
rect 4904 -10898 4938 -9946
rect 5288 -10898 5322 -9946
rect 5824 -10898 5858 -9946
rect 1709 -10994 2077 -10960
rect 2629 -10994 2997 -10960
rect 3549 -10994 3917 -10960
rect 4469 -10994 4837 -10960
rect 5389 -10994 5757 -10960
rect 6392 -10164 6560 -10130
rect 6330 -10299 6364 -10223
rect 6588 -10299 6622 -10223
rect 6670 -10320 6702 -10200
rect 6702 -10320 6736 -10200
rect 6736 -10320 6760 -10200
rect 6392 -10392 6560 -10358
rect 6392 -10732 6560 -10698
rect 6330 -10858 6364 -10782
rect 6588 -10858 6622 -10782
rect 6392 -10942 6560 -10908
<< metal1 >>
rect -1386 2642 -1136 2650
rect 284 2642 674 2650
rect -1386 2626 2093 2642
rect -1386 2592 -1127 2626
rect -1093 2592 -1029 2626
rect -995 2592 -931 2626
rect -897 2592 -833 2626
rect -799 2592 -735 2626
rect -701 2592 -637 2626
rect -603 2592 -539 2626
rect -505 2592 -441 2626
rect -407 2592 -343 2626
rect -309 2592 -245 2626
rect -211 2592 -147 2626
rect -113 2592 -49 2626
rect -15 2592 49 2626
rect 83 2592 147 2626
rect 181 2592 245 2626
rect 279 2592 671 2626
rect 705 2592 769 2626
rect 803 2592 867 2626
rect 901 2592 965 2626
rect 999 2592 1063 2626
rect 1097 2592 1161 2626
rect 1195 2592 1259 2626
rect 1293 2592 1357 2626
rect 1391 2592 1455 2626
rect 1489 2592 1553 2626
rect 1587 2592 1651 2626
rect 1685 2592 1749 2626
rect 1783 2592 1847 2626
rect 1881 2592 1945 2626
rect 1979 2592 2043 2626
rect 2077 2592 2093 2626
rect -1386 2580 2093 2592
rect -1386 2110 -1236 2580
rect -1143 2576 295 2580
rect -1182 2533 -1136 2545
rect -1182 2305 -1176 2533
rect -1142 2305 -1136 2533
rect -1097 2385 -1087 2545
rect -1035 2385 -1025 2545
rect -986 2533 -940 2545
rect -1195 2145 -1185 2305
rect -1133 2145 -1123 2305
rect -1084 2157 -1078 2385
rect -1044 2157 -1038 2385
rect -986 2305 -980 2533
rect -946 2305 -940 2533
rect -901 2385 -891 2545
rect -839 2385 -829 2545
rect -790 2533 -744 2545
rect -1084 2145 -1038 2157
rect -999 2145 -989 2305
rect -937 2145 -927 2305
rect -888 2157 -882 2385
rect -848 2157 -842 2385
rect -790 2305 -784 2533
rect -750 2305 -744 2533
rect -705 2385 -695 2545
rect -643 2385 -633 2545
rect -594 2533 -548 2545
rect -888 2145 -842 2157
rect -803 2145 -793 2305
rect -741 2145 -731 2305
rect -692 2157 -686 2385
rect -652 2157 -646 2385
rect -594 2305 -588 2533
rect -554 2305 -548 2533
rect -509 2385 -499 2545
rect -447 2385 -437 2545
rect -398 2533 -352 2545
rect -692 2145 -646 2157
rect -607 2145 -597 2305
rect -545 2145 -535 2305
rect -496 2157 -490 2385
rect -456 2157 -450 2385
rect -398 2305 -392 2533
rect -358 2305 -352 2533
rect -313 2385 -303 2545
rect -251 2385 -241 2545
rect -202 2533 -156 2545
rect -496 2145 -450 2157
rect -411 2145 -401 2305
rect -349 2145 -339 2305
rect -300 2157 -294 2385
rect -260 2157 -254 2385
rect -202 2305 -196 2533
rect -162 2305 -156 2533
rect -117 2385 -107 2545
rect -55 2385 -45 2545
rect -6 2533 40 2545
rect -300 2145 -254 2157
rect -215 2145 -205 2305
rect -153 2145 -143 2305
rect -104 2157 -98 2385
rect -64 2157 -58 2385
rect -6 2305 0 2533
rect 34 2305 40 2533
rect 79 2385 89 2545
rect 141 2385 151 2545
rect 190 2533 236 2545
rect -104 2145 -58 2157
rect -19 2145 -9 2305
rect 43 2145 53 2305
rect 92 2157 98 2385
rect 132 2157 138 2385
rect 190 2305 196 2533
rect 230 2305 236 2533
rect 275 2385 285 2545
rect 337 2385 347 2545
rect 92 2145 138 2157
rect 177 2145 187 2305
rect 239 2145 249 2305
rect 288 2157 294 2385
rect 328 2157 334 2385
rect 288 2145 334 2157
rect -1143 2110 295 2114
rect 434 2110 514 2580
rect 655 2576 2093 2580
rect 616 2533 662 2545
rect 616 2305 622 2533
rect 656 2305 662 2533
rect 701 2385 711 2545
rect 763 2385 773 2545
rect 812 2533 858 2545
rect 603 2145 613 2305
rect 665 2145 675 2305
rect 714 2157 720 2385
rect 754 2157 760 2385
rect 812 2305 818 2533
rect 852 2305 858 2533
rect 897 2385 907 2545
rect 959 2385 969 2545
rect 1008 2533 1054 2545
rect 714 2145 760 2157
rect 799 2145 809 2305
rect 861 2145 871 2305
rect 910 2157 916 2385
rect 950 2157 956 2385
rect 1008 2305 1014 2533
rect 1048 2305 1054 2533
rect 1093 2385 1103 2545
rect 1155 2385 1165 2545
rect 1204 2533 1250 2545
rect 910 2145 956 2157
rect 995 2145 1005 2305
rect 1057 2145 1067 2305
rect 1106 2157 1112 2385
rect 1146 2157 1152 2385
rect 1204 2305 1210 2533
rect 1244 2305 1250 2533
rect 1289 2385 1299 2545
rect 1351 2385 1361 2545
rect 1400 2533 1446 2545
rect 1106 2145 1152 2157
rect 1191 2145 1201 2305
rect 1253 2145 1263 2305
rect 1302 2157 1308 2385
rect 1342 2157 1348 2385
rect 1400 2305 1406 2533
rect 1440 2305 1446 2533
rect 1485 2385 1495 2545
rect 1547 2385 1557 2545
rect 1596 2533 1642 2545
rect 1302 2145 1348 2157
rect 1387 2145 1397 2305
rect 1449 2145 1459 2305
rect 1498 2157 1504 2385
rect 1538 2157 1544 2385
rect 1596 2305 1602 2533
rect 1636 2305 1642 2533
rect 1681 2385 1691 2545
rect 1743 2385 1753 2545
rect 1792 2533 1838 2545
rect 1498 2145 1544 2157
rect 1583 2145 1593 2305
rect 1645 2145 1655 2305
rect 1694 2157 1700 2385
rect 1734 2157 1740 2385
rect 1792 2305 1798 2533
rect 1832 2305 1838 2533
rect 1877 2385 1887 2545
rect 1939 2385 1949 2545
rect 1988 2533 2034 2545
rect 1694 2145 1740 2157
rect 1779 2145 1789 2305
rect 1841 2145 1851 2305
rect 1890 2157 1896 2385
rect 1930 2157 1936 2385
rect 1988 2305 1994 2533
rect 2028 2305 2034 2533
rect 2073 2385 2083 2545
rect 2135 2385 2145 2545
rect 1890 2145 1936 2157
rect 1975 2145 1985 2305
rect 2037 2145 2047 2305
rect 2086 2157 2092 2385
rect 2126 2157 2132 2385
rect 2086 2145 2132 2157
rect 655 2110 2093 2114
rect -1386 2098 2104 2110
rect -1386 2064 -1127 2098
rect -1093 2064 -1029 2098
rect -995 2064 -931 2098
rect -897 2064 -833 2098
rect -799 2064 -735 2098
rect -701 2064 -637 2098
rect -603 2064 -539 2098
rect -505 2064 -441 2098
rect -407 2064 -343 2098
rect -309 2064 -245 2098
rect -211 2064 -147 2098
rect -113 2064 -49 2098
rect -15 2064 49 2098
rect 83 2064 147 2098
rect 181 2064 245 2098
rect 279 2064 671 2098
rect 705 2064 769 2098
rect 803 2064 867 2098
rect 901 2064 965 2098
rect 999 2064 1063 2098
rect 1097 2064 1161 2098
rect 1195 2064 1259 2098
rect 1293 2064 1357 2098
rect 1391 2064 1455 2098
rect 1489 2064 1553 2098
rect 1587 2064 1651 2098
rect 1685 2064 1749 2098
rect 1783 2064 1847 2098
rect 1881 2064 1945 2098
rect 1979 2064 2043 2098
rect 2077 2064 2104 2098
rect 2208 2070 2350 2082
rect -1386 1990 2104 2064
rect -1386 1956 -1127 1990
rect -1093 1956 -1029 1990
rect -995 1956 -931 1990
rect -897 1956 -833 1990
rect -799 1956 -735 1990
rect -701 1956 -637 1990
rect -603 1956 -539 1990
rect -505 1956 -441 1990
rect -407 1956 -343 1990
rect -309 1956 -245 1990
rect -211 1956 -147 1990
rect -113 1956 -49 1990
rect -15 1956 49 1990
rect 83 1956 147 1990
rect 181 1956 245 1990
rect 279 1956 671 1990
rect 705 1956 769 1990
rect 803 1956 867 1990
rect 901 1956 965 1990
rect 999 1956 1063 1990
rect 1097 1956 1161 1990
rect 1195 1956 1259 1990
rect 1293 1956 1357 1990
rect 1391 1956 1455 1990
rect 1489 1956 1553 1990
rect 1587 1956 1651 1990
rect 1685 1956 1749 1990
rect 1783 1956 1847 1990
rect 1881 1956 1945 1990
rect 1979 1956 2043 1990
rect 2077 1956 2104 1990
rect -1386 1940 2104 1956
rect -1386 1470 -1236 1940
rect -1195 1749 -1185 1909
rect -1133 1749 -1123 1909
rect -1084 1897 -1038 1909
rect -1182 1521 -1176 1749
rect -1142 1521 -1136 1749
rect -1084 1669 -1078 1897
rect -1044 1669 -1038 1897
rect -999 1749 -989 1909
rect -937 1749 -927 1909
rect -888 1897 -842 1909
rect -1182 1509 -1136 1521
rect -1097 1509 -1087 1669
rect -1035 1509 -1025 1669
rect -986 1521 -980 1749
rect -946 1521 -940 1749
rect -888 1669 -882 1897
rect -848 1669 -842 1897
rect -803 1749 -793 1909
rect -741 1749 -731 1909
rect -692 1897 -646 1909
rect -986 1509 -940 1521
rect -901 1509 -891 1669
rect -839 1509 -829 1669
rect -790 1521 -784 1749
rect -750 1521 -744 1749
rect -692 1669 -686 1897
rect -652 1669 -646 1897
rect -607 1749 -597 1909
rect -545 1749 -535 1909
rect -496 1897 -450 1909
rect -790 1509 -744 1521
rect -705 1509 -695 1669
rect -643 1509 -633 1669
rect -594 1521 -588 1749
rect -554 1521 -548 1749
rect -496 1669 -490 1897
rect -456 1669 -450 1897
rect -411 1749 -401 1909
rect -349 1749 -339 1909
rect -300 1897 -254 1909
rect -594 1509 -548 1521
rect -509 1509 -499 1669
rect -447 1509 -437 1669
rect -398 1521 -392 1749
rect -358 1521 -352 1749
rect -300 1669 -294 1897
rect -260 1669 -254 1897
rect -215 1749 -205 1909
rect -153 1749 -143 1909
rect -104 1897 -58 1909
rect -398 1509 -352 1521
rect -313 1509 -303 1669
rect -251 1509 -241 1669
rect -202 1521 -196 1749
rect -162 1521 -156 1749
rect -104 1669 -98 1897
rect -64 1669 -58 1897
rect -19 1749 -9 1909
rect 43 1749 53 1909
rect 92 1897 138 1909
rect -202 1509 -156 1521
rect -117 1509 -107 1669
rect -55 1509 -45 1669
rect -6 1521 0 1749
rect 34 1521 40 1749
rect 92 1669 98 1897
rect 132 1669 138 1897
rect 177 1749 187 1909
rect 239 1749 249 1909
rect 288 1897 334 1909
rect -6 1509 40 1521
rect 79 1509 89 1669
rect 141 1509 151 1669
rect 190 1521 196 1749
rect 230 1521 236 1749
rect 288 1669 294 1897
rect 328 1669 334 1897
rect 190 1509 236 1521
rect 275 1509 285 1669
rect 337 1509 347 1669
rect 434 1480 514 1940
rect 603 1749 613 1909
rect 665 1749 675 1909
rect 714 1897 760 1909
rect 616 1521 622 1749
rect 656 1521 662 1749
rect 714 1669 720 1897
rect 754 1669 760 1897
rect 799 1749 809 1909
rect 861 1749 871 1909
rect 910 1897 956 1909
rect 616 1509 662 1521
rect 701 1509 711 1669
rect 763 1509 773 1669
rect 812 1521 818 1749
rect 852 1521 858 1749
rect 910 1669 916 1897
rect 950 1669 956 1897
rect 995 1749 1005 1909
rect 1057 1749 1067 1909
rect 1106 1897 1152 1909
rect 812 1509 858 1521
rect 897 1509 907 1669
rect 959 1509 969 1669
rect 1008 1521 1014 1749
rect 1048 1521 1054 1749
rect 1106 1669 1112 1897
rect 1146 1669 1152 1897
rect 1191 1749 1201 1909
rect 1253 1749 1263 1909
rect 1302 1897 1348 1909
rect 1008 1509 1054 1521
rect 1093 1509 1103 1669
rect 1155 1509 1165 1669
rect 1204 1521 1210 1749
rect 1244 1521 1250 1749
rect 1302 1669 1308 1897
rect 1342 1669 1348 1897
rect 1387 1749 1397 1909
rect 1449 1749 1459 1909
rect 1498 1897 1544 1909
rect 1204 1509 1250 1521
rect 1289 1509 1299 1669
rect 1351 1509 1361 1669
rect 1400 1521 1406 1749
rect 1440 1521 1446 1749
rect 1498 1669 1504 1897
rect 1538 1669 1544 1897
rect 1583 1749 1593 1909
rect 1645 1749 1655 1909
rect 1694 1897 1740 1909
rect 1400 1509 1446 1521
rect 1485 1509 1495 1669
rect 1547 1509 1557 1669
rect 1596 1521 1602 1749
rect 1636 1521 1642 1749
rect 1694 1669 1700 1897
rect 1734 1669 1740 1897
rect 1779 1749 1789 1909
rect 1841 1749 1851 1909
rect 1890 1897 1936 1909
rect 1596 1509 1642 1521
rect 1681 1509 1691 1669
rect 1743 1509 1753 1669
rect 1792 1521 1798 1749
rect 1832 1521 1838 1749
rect 1890 1669 1896 1897
rect 1930 1669 1936 1897
rect 1975 1749 1985 1909
rect 2037 1749 2047 1909
rect 2086 1897 2132 1909
rect 1792 1509 1838 1521
rect 1877 1509 1887 1669
rect 1939 1509 1949 1669
rect 1988 1521 1994 1749
rect 2028 1521 2034 1749
rect 2086 1669 2092 1897
rect 2126 1669 2132 1897
rect 1988 1509 2034 1521
rect 2073 1509 2083 1669
rect 2135 1509 2145 1669
rect 2204 1510 2214 2070
rect 2344 1510 2354 2070
rect 4100 1996 4660 2000
rect 4098 1980 4660 1996
rect 2474 1974 4660 1980
rect 2474 1940 2486 1974
rect 2554 1940 2644 1974
rect 2712 1940 2802 1974
rect 2870 1940 2960 1974
rect 3028 1940 3118 1974
rect 3186 1940 3276 1974
rect 3344 1940 3434 1974
rect 3502 1940 3592 1974
rect 3660 1940 3750 1974
rect 3818 1940 3908 1974
rect 3976 1940 4660 1974
rect 2474 1934 2566 1940
rect 2632 1934 2724 1940
rect 2790 1934 2882 1940
rect 2948 1934 3040 1940
rect 3106 1934 3198 1940
rect 3264 1934 3356 1940
rect 3422 1934 3514 1940
rect 3580 1934 3672 1940
rect 3738 1934 3830 1940
rect 3896 1934 3988 1940
rect 4094 1930 4660 1940
rect 4740 1930 4750 2000
rect 2418 1881 2464 1893
rect 2418 1653 2424 1881
rect 2458 1653 2464 1881
rect 2563 1733 2573 1893
rect 2625 1733 2635 1893
rect 2734 1881 2780 1893
rect 2208 1498 2350 1510
rect 2405 1493 2415 1653
rect 2467 1493 2477 1653
rect 2576 1505 2582 1733
rect 2616 1505 2622 1733
rect 2734 1653 2740 1881
rect 2774 1653 2780 1881
rect 2879 1733 2889 1893
rect 2941 1733 2951 1893
rect 3050 1881 3096 1893
rect 2576 1493 2622 1505
rect 2721 1493 2731 1653
rect 2783 1493 2793 1653
rect 2892 1505 2898 1733
rect 2932 1505 2938 1733
rect 3050 1653 3056 1881
rect 3090 1653 3096 1881
rect 3195 1733 3205 1893
rect 3257 1733 3267 1893
rect 3366 1881 3412 1893
rect 2892 1493 2938 1505
rect 3037 1493 3047 1653
rect 3099 1493 3109 1653
rect 3208 1505 3214 1733
rect 3248 1505 3254 1733
rect 3366 1653 3372 1881
rect 3406 1653 3412 1881
rect 3511 1733 3521 1893
rect 3573 1733 3583 1893
rect 3682 1881 3728 1893
rect 3208 1493 3254 1505
rect 3353 1493 3363 1653
rect 3415 1493 3425 1653
rect 3524 1505 3530 1733
rect 3564 1505 3570 1733
rect 3682 1653 3688 1881
rect 3722 1653 3728 1881
rect 3827 1733 3837 1893
rect 3889 1733 3899 1893
rect 3998 1881 4044 1893
rect 3524 1493 3570 1505
rect 3669 1493 3679 1653
rect 3731 1493 3741 1653
rect 3840 1505 3846 1733
rect 3880 1505 3886 1733
rect 3998 1653 4004 1881
rect 4038 1653 4044 1881
rect 3840 1493 3886 1505
rect 3985 1493 3995 1653
rect 4047 1493 4057 1653
rect 284 1478 674 1480
rect -1143 1470 2093 1478
rect -1386 1462 2093 1470
rect -1386 1428 -1127 1462
rect -1093 1428 -1029 1462
rect -995 1428 -931 1462
rect -897 1428 -833 1462
rect -799 1428 -735 1462
rect -701 1428 -637 1462
rect -603 1428 -539 1462
rect -505 1428 -441 1462
rect -407 1428 -343 1462
rect -309 1428 -245 1462
rect -211 1428 -147 1462
rect -113 1428 -49 1462
rect -15 1428 49 1462
rect 83 1428 147 1462
rect 181 1428 245 1462
rect 279 1428 671 1462
rect 705 1428 769 1462
rect 803 1428 867 1462
rect 901 1428 965 1462
rect 999 1428 1063 1462
rect 1097 1428 1161 1462
rect 1195 1428 1259 1462
rect 1293 1428 1357 1462
rect 1391 1428 1455 1462
rect 1489 1428 1553 1462
rect 1587 1428 1651 1462
rect 1685 1428 1749 1462
rect 1783 1428 1847 1462
rect 1881 1428 1945 1462
rect 1979 1428 2043 1462
rect 2077 1428 2093 1462
rect 2474 1446 2566 1452
rect 2474 1440 2486 1446
rect -1386 1412 2093 1428
rect 2464 1412 2486 1440
rect 2554 1440 2566 1446
rect 2632 1446 2724 1452
rect 2632 1440 2644 1446
rect 2554 1412 2644 1440
rect 2712 1440 2724 1446
rect 2790 1446 2882 1452
rect 2790 1440 2802 1446
rect 2712 1412 2802 1440
rect 2870 1440 2882 1446
rect 2948 1446 3040 1452
rect 2948 1440 2960 1446
rect 2870 1412 2960 1440
rect 3028 1440 3040 1446
rect 3106 1446 3198 1452
rect 3106 1440 3118 1446
rect 3028 1412 3118 1440
rect 3186 1440 3198 1446
rect 3264 1446 3356 1452
rect 3264 1440 3276 1446
rect 3186 1412 3276 1440
rect 3344 1440 3356 1446
rect 3422 1446 3514 1452
rect 3422 1440 3434 1446
rect 3344 1412 3434 1440
rect 3502 1440 3514 1446
rect 3580 1446 3672 1452
rect 3580 1440 3592 1446
rect 3502 1412 3592 1440
rect 3660 1440 3672 1446
rect 3738 1446 3830 1452
rect 3738 1440 3750 1446
rect 3660 1412 3750 1440
rect 3818 1440 3830 1446
rect 3896 1446 3988 1452
rect 3896 1440 3908 1446
rect 3818 1412 3908 1440
rect 3976 1440 3988 1446
rect 4094 1440 4134 1930
rect 3976 1412 4134 1440
rect -1386 1400 -1136 1412
rect 284 1410 674 1412
rect -1386 1180 -1236 1400
rect 434 1220 514 1410
rect 2464 1400 4134 1412
rect -1386 1166 -1136 1180
rect 434 1166 1544 1220
rect -1386 1150 1544 1166
rect -1386 1116 -1127 1150
rect -1093 1116 -1030 1150
rect -996 1116 -931 1150
rect -897 1116 -834 1150
rect -800 1116 -735 1150
rect -701 1116 -638 1150
rect -604 1116 -539 1150
rect -505 1116 -442 1150
rect -408 1116 -343 1150
rect -309 1116 -246 1150
rect -212 1116 -147 1150
rect -113 1116 -50 1150
rect -16 1116 49 1150
rect 83 1116 146 1150
rect 180 1116 245 1150
rect 279 1116 342 1150
rect 376 1116 441 1150
rect 475 1116 538 1150
rect 572 1116 637 1150
rect 671 1116 734 1150
rect 768 1116 833 1150
rect 867 1116 930 1150
rect 964 1116 1029 1150
rect 1063 1116 1126 1150
rect 1160 1116 1225 1150
rect 1259 1116 1544 1150
rect -1386 1110 1544 1116
rect -1386 640 -1236 1110
rect -1144 1106 1274 1110
rect -1182 1066 -1136 1078
rect -1182 838 -1176 1066
rect -1142 838 -1136 1066
rect -1097 918 -1087 1078
rect -1035 918 -1025 1078
rect -986 1066 -940 1078
rect -1195 678 -1185 838
rect -1133 678 -1123 838
rect -1084 690 -1078 918
rect -1044 690 -1038 918
rect -986 838 -980 1066
rect -946 838 -940 1066
rect -901 918 -891 1078
rect -839 918 -829 1078
rect -790 1066 -744 1078
rect -1084 678 -1038 690
rect -999 678 -989 838
rect -937 678 -927 838
rect -888 690 -882 918
rect -848 690 -842 918
rect -790 838 -784 1066
rect -750 838 -744 1066
rect -705 918 -695 1078
rect -643 918 -633 1078
rect -594 1066 -548 1078
rect -888 678 -842 690
rect -803 678 -793 838
rect -741 678 -731 838
rect -692 690 -686 918
rect -652 690 -646 918
rect -594 838 -588 1066
rect -554 838 -548 1066
rect -509 918 -499 1078
rect -447 918 -437 1078
rect -398 1066 -352 1078
rect -692 678 -646 690
rect -607 678 -597 838
rect -545 678 -535 838
rect -496 690 -490 918
rect -456 690 -450 918
rect -398 838 -392 1066
rect -358 838 -352 1066
rect -313 918 -303 1078
rect -251 918 -241 1078
rect -202 1066 -156 1078
rect -496 678 -450 690
rect -411 678 -401 838
rect -349 678 -339 838
rect -300 690 -294 918
rect -260 690 -254 918
rect -202 838 -196 1066
rect -162 838 -156 1066
rect -117 918 -107 1078
rect -55 918 -45 1078
rect -6 1066 40 1078
rect -300 678 -254 690
rect -215 678 -205 838
rect -153 678 -143 838
rect -104 690 -98 918
rect -64 690 -58 918
rect -6 838 0 1066
rect 34 838 40 1066
rect 79 918 89 1078
rect 141 918 151 1078
rect 190 1066 236 1078
rect -104 678 -58 690
rect -19 678 -9 838
rect 43 678 53 838
rect 92 690 98 918
rect 132 690 138 918
rect 190 838 196 1066
rect 230 838 236 1066
rect 275 918 285 1078
rect 337 918 347 1078
rect 386 1066 432 1078
rect 92 678 138 690
rect 177 678 187 838
rect 239 678 249 838
rect 288 690 294 918
rect 328 690 334 918
rect 386 838 392 1066
rect 426 838 432 1066
rect 471 918 481 1078
rect 533 918 543 1078
rect 582 1066 628 1078
rect 288 678 334 690
rect 373 678 383 838
rect 435 678 445 838
rect 484 690 490 918
rect 524 690 530 918
rect 582 838 588 1066
rect 622 838 628 1066
rect 667 918 677 1078
rect 729 918 739 1078
rect 778 1066 824 1078
rect 484 678 530 690
rect 569 678 579 838
rect 631 678 641 838
rect 680 690 686 918
rect 720 690 726 918
rect 778 838 784 1066
rect 818 838 824 1066
rect 863 918 873 1078
rect 925 918 935 1078
rect 974 1066 1020 1078
rect 680 678 726 690
rect 765 678 775 838
rect 827 678 837 838
rect 876 690 882 918
rect 916 690 922 918
rect 974 838 980 1066
rect 1014 838 1020 1066
rect 1059 918 1069 1078
rect 1121 918 1131 1078
rect 1170 1066 1216 1078
rect 876 678 922 690
rect 961 678 971 838
rect 1023 678 1033 838
rect 1072 690 1078 918
rect 1112 690 1118 918
rect 1170 838 1176 1066
rect 1210 838 1216 1066
rect 1255 918 1265 1078
rect 1317 918 1327 1078
rect 1072 678 1118 690
rect 1157 678 1167 838
rect 1219 678 1229 838
rect 1268 690 1274 918
rect 1308 690 1314 918
rect 1268 678 1314 690
rect -1144 640 1274 650
rect 1404 640 1544 1110
rect 2154 660 2164 850
rect 2414 846 3954 850
rect 2414 830 3955 846
rect 2414 796 2533 830
rect 2567 796 2631 830
rect 2665 796 2729 830
rect 2763 796 2827 830
rect 2861 796 2925 830
rect 2959 796 3023 830
rect 3057 796 3121 830
rect 3155 796 3219 830
rect 3253 796 3317 830
rect 3351 796 3415 830
rect 3449 796 3513 830
rect 3547 796 3611 830
rect 3645 796 3709 830
rect 3743 796 3807 830
rect 3841 796 3905 830
rect 3939 796 3955 830
rect 2414 790 3955 796
rect 2414 660 2434 790
rect -1386 606 -1128 640
rect -1094 606 -1029 640
rect -995 606 -932 640
rect -898 606 -833 640
rect -799 606 -736 640
rect -702 606 -637 640
rect -603 606 -540 640
rect -506 606 -441 640
rect -407 606 -344 640
rect -310 606 -245 640
rect -211 606 -148 640
rect -114 606 -49 640
rect -15 606 48 640
rect 82 606 147 640
rect 181 606 244 640
rect 278 606 343 640
rect 377 606 440 640
rect 474 606 539 640
rect 573 606 636 640
rect 670 606 735 640
rect 769 606 832 640
rect 866 606 931 640
rect 965 606 1028 640
rect 1062 606 1127 640
rect 1161 606 1224 640
rect 1258 606 1544 640
rect -1386 532 1544 606
rect -1386 498 -1127 532
rect -1093 498 -1029 532
rect -995 498 -931 532
rect -897 498 -833 532
rect -799 498 -735 532
rect -701 498 -637 532
rect -603 498 -539 532
rect -505 498 -441 532
rect -407 498 -343 532
rect -309 498 -245 532
rect -211 498 -147 532
rect -113 498 -49 532
rect -15 498 49 532
rect 83 498 147 532
rect 181 498 245 532
rect 279 498 343 532
rect 377 498 441 532
rect 475 498 539 532
rect 573 498 637 532
rect 671 498 735 532
rect 769 498 833 532
rect 867 498 931 532
rect 965 498 1029 532
rect 1063 498 1127 532
rect 1161 498 1225 532
rect 1259 498 1544 532
rect -1386 490 1544 498
rect -1386 30 -1236 490
rect -1143 488 1275 490
rect -1195 300 -1185 460
rect -1133 300 -1123 460
rect -1084 448 -1038 460
rect -1182 72 -1176 300
rect -1142 72 -1136 300
rect -1084 220 -1078 448
rect -1044 220 -1038 448
rect -999 300 -989 460
rect -937 300 -927 460
rect -888 448 -842 460
rect -1182 60 -1136 72
rect -1097 60 -1087 220
rect -1035 60 -1025 220
rect -986 72 -980 300
rect -946 72 -940 300
rect -888 220 -882 448
rect -848 220 -842 448
rect -803 300 -793 460
rect -741 300 -731 460
rect -692 448 -646 460
rect -986 60 -940 72
rect -901 60 -891 220
rect -839 60 -829 220
rect -790 72 -784 300
rect -750 72 -744 300
rect -692 220 -686 448
rect -652 220 -646 448
rect -607 300 -597 460
rect -545 300 -535 460
rect -496 448 -450 460
rect -790 60 -744 72
rect -705 60 -695 220
rect -643 60 -633 220
rect -594 72 -588 300
rect -554 72 -548 300
rect -496 220 -490 448
rect -456 220 -450 448
rect -411 300 -401 460
rect -349 300 -339 460
rect -300 448 -254 460
rect -594 60 -548 72
rect -509 60 -499 220
rect -447 60 -437 220
rect -398 72 -392 300
rect -358 72 -352 300
rect -300 220 -294 448
rect -260 220 -254 448
rect -215 300 -205 460
rect -153 300 -143 460
rect -104 448 -58 460
rect -398 60 -352 72
rect -313 60 -303 220
rect -251 60 -241 220
rect -202 72 -196 300
rect -162 72 -156 300
rect -104 220 -98 448
rect -64 220 -58 448
rect -19 300 -9 460
rect 43 300 53 460
rect 92 448 138 460
rect -202 60 -156 72
rect -117 60 -107 220
rect -55 60 -45 220
rect -6 72 0 300
rect 34 72 40 300
rect 92 220 98 448
rect 132 220 138 448
rect 177 300 187 460
rect 239 300 249 460
rect 288 448 334 460
rect -6 60 40 72
rect 79 60 89 220
rect 141 60 151 220
rect 190 72 196 300
rect 230 72 236 300
rect 288 220 294 448
rect 328 220 334 448
rect 373 300 383 460
rect 435 300 445 460
rect 484 448 530 460
rect 190 60 236 72
rect 275 60 285 220
rect 337 60 347 220
rect 386 72 392 300
rect 426 72 432 300
rect 484 220 490 448
rect 524 220 530 448
rect 569 300 579 460
rect 631 300 641 460
rect 680 448 726 460
rect 386 60 432 72
rect 471 60 481 220
rect 533 60 543 220
rect 582 72 588 300
rect 622 72 628 300
rect 680 220 686 448
rect 720 220 726 448
rect 765 300 775 460
rect 827 300 837 460
rect 876 448 922 460
rect 582 60 628 72
rect 667 60 677 220
rect 729 60 739 220
rect 778 72 784 300
rect 818 72 824 300
rect 876 220 882 448
rect 916 220 922 448
rect 961 300 971 460
rect 1023 300 1033 460
rect 1072 448 1118 460
rect 778 60 824 72
rect 863 60 873 220
rect 925 60 935 220
rect 974 72 980 300
rect 1014 72 1020 300
rect 1072 220 1078 448
rect 1112 220 1118 448
rect 1157 300 1167 460
rect 1219 300 1229 460
rect 1268 448 1314 460
rect 974 60 1020 72
rect 1059 60 1069 220
rect 1121 60 1131 220
rect 1170 72 1176 300
rect 1210 72 1216 300
rect 1268 220 1274 448
rect 1308 220 1314 448
rect 1404 320 1544 490
rect 2198 320 2290 332
rect 2344 320 2434 660
rect 2465 598 2475 758
rect 2527 598 2537 758
rect 2576 746 2622 758
rect 2478 370 2484 598
rect 2518 370 2524 598
rect 2576 518 2582 746
rect 2616 518 2622 746
rect 2661 598 2671 758
rect 2723 598 2733 758
rect 2772 746 2818 758
rect 2478 358 2524 370
rect 2563 358 2573 518
rect 2625 358 2635 518
rect 2674 370 2680 598
rect 2714 370 2720 598
rect 2772 518 2778 746
rect 2812 518 2818 746
rect 2857 598 2867 758
rect 2919 598 2929 758
rect 2968 746 3014 758
rect 2674 358 2720 370
rect 2759 358 2769 518
rect 2821 358 2831 518
rect 2870 370 2876 598
rect 2910 370 2916 598
rect 2968 518 2974 746
rect 3008 518 3014 746
rect 3053 598 3063 758
rect 3115 598 3125 758
rect 3164 746 3210 758
rect 2870 358 2916 370
rect 2955 358 2965 518
rect 3017 358 3027 518
rect 3066 370 3072 598
rect 3106 370 3112 598
rect 3164 518 3170 746
rect 3204 518 3210 746
rect 3249 598 3259 758
rect 3311 598 3321 758
rect 3360 746 3406 758
rect 3066 358 3112 370
rect 3151 358 3161 518
rect 3213 358 3223 518
rect 3262 370 3268 598
rect 3302 370 3308 598
rect 3360 518 3366 746
rect 3400 518 3406 746
rect 3445 598 3455 758
rect 3507 598 3517 758
rect 3556 746 3602 758
rect 3262 358 3308 370
rect 3347 358 3357 518
rect 3409 358 3419 518
rect 3458 370 3464 598
rect 3498 370 3504 598
rect 3556 518 3562 746
rect 3596 518 3602 746
rect 3641 598 3651 758
rect 3703 598 3713 758
rect 3752 746 3798 758
rect 3458 358 3504 370
rect 3543 358 3553 518
rect 3605 358 3615 518
rect 3654 370 3660 598
rect 3694 370 3700 598
rect 3752 518 3758 746
rect 3792 518 3798 746
rect 3837 598 3847 758
rect 3899 598 3909 758
rect 3948 746 3994 758
rect 3654 358 3700 370
rect 3739 358 3749 518
rect 3801 358 3811 518
rect 3850 370 3856 598
rect 3890 370 3896 598
rect 3948 518 3954 746
rect 3988 518 3994 746
rect 3850 358 3896 370
rect 3935 358 3945 518
rect 3997 358 4007 518
rect 4048 340 4180 352
rect 2517 320 3955 326
rect 1170 60 1216 72
rect 1255 60 1265 220
rect 1317 60 1327 220
rect 1404 160 1454 320
rect 1684 160 1694 320
rect 2194 160 2204 320
rect 2284 160 2294 320
rect 2344 286 2533 320
rect 2567 286 2631 320
rect 2665 286 2729 320
rect 2763 286 2827 320
rect 2861 286 2925 320
rect 2959 286 3023 320
rect 3057 286 3121 320
rect 3155 286 3219 320
rect 3253 286 3317 320
rect 3351 286 3415 320
rect 3449 286 3513 320
rect 3547 286 3611 320
rect 3645 286 3709 320
rect 3743 286 3807 320
rect 3841 286 3905 320
rect 3939 286 3955 320
rect 2344 270 3955 286
rect 2344 228 3954 270
rect 2344 212 3955 228
rect 2344 180 2533 212
rect -1143 30 1275 32
rect 1404 30 1544 160
rect 2198 148 2290 160
rect -1386 22 1544 30
rect -1386 -12 -1127 22
rect -1093 -12 -1029 22
rect -995 -12 -931 22
rect -897 -12 -833 22
rect -799 -12 -735 22
rect -701 -12 -637 22
rect -603 -12 -539 22
rect -505 -12 -441 22
rect -407 -12 -343 22
rect -309 -12 -245 22
rect -211 -12 -147 22
rect -113 -12 -49 22
rect -15 -12 49 22
rect 83 -12 147 22
rect 181 -12 245 22
rect 279 -12 343 22
rect 377 -12 441 22
rect 475 -12 539 22
rect 573 -12 637 22
rect 671 -12 735 22
rect 769 -12 833 22
rect 867 -12 931 22
rect 965 -12 1029 22
rect 1063 -12 1127 22
rect 1161 -12 1225 22
rect 1259 -12 1544 22
rect -1386 -28 1544 -12
rect -1386 -30 -1136 -28
rect 1274 -30 1544 -28
rect -1386 -260 -1236 -30
rect -1386 -278 -1136 -260
rect 1404 -270 1544 -30
rect 1274 -278 1544 -270
rect -1386 -294 1544 -278
rect -1386 -328 -1127 -294
rect -1093 -328 -1030 -294
rect -996 -328 -931 -294
rect -897 -328 -834 -294
rect -800 -328 -735 -294
rect -701 -328 -638 -294
rect -604 -328 -539 -294
rect -505 -328 -442 -294
rect -408 -328 -343 -294
rect -309 -328 -246 -294
rect -212 -328 -147 -294
rect -113 -328 -50 -294
rect -16 -328 49 -294
rect 83 -328 146 -294
rect 180 -328 245 -294
rect 279 -328 342 -294
rect 376 -328 441 -294
rect 475 -328 538 -294
rect 572 -328 637 -294
rect 671 -328 734 -294
rect 768 -328 833 -294
rect 867 -328 930 -294
rect 964 -328 1029 -294
rect 1063 -328 1126 -294
rect 1160 -328 1225 -294
rect 1259 -328 1544 -294
rect -1386 -330 1544 -328
rect -1386 -800 -1236 -330
rect -1144 -338 1274 -330
rect -1182 -378 -1136 -366
rect -1182 -606 -1176 -378
rect -1142 -606 -1136 -378
rect -1097 -526 -1087 -366
rect -1035 -526 -1025 -366
rect -986 -378 -940 -366
rect -1195 -766 -1185 -606
rect -1133 -766 -1123 -606
rect -1084 -754 -1078 -526
rect -1044 -754 -1038 -526
rect -986 -606 -980 -378
rect -946 -606 -940 -378
rect -901 -526 -891 -366
rect -839 -526 -829 -366
rect -790 -378 -744 -366
rect -1084 -766 -1038 -754
rect -999 -766 -989 -606
rect -937 -766 -927 -606
rect -888 -754 -882 -526
rect -848 -754 -842 -526
rect -790 -606 -784 -378
rect -750 -606 -744 -378
rect -705 -526 -695 -366
rect -643 -526 -633 -366
rect -594 -378 -548 -366
rect -888 -766 -842 -754
rect -803 -766 -793 -606
rect -741 -766 -731 -606
rect -692 -754 -686 -526
rect -652 -754 -646 -526
rect -594 -606 -588 -378
rect -554 -606 -548 -378
rect -509 -526 -499 -366
rect -447 -526 -437 -366
rect -398 -378 -352 -366
rect -692 -766 -646 -754
rect -607 -766 -597 -606
rect -545 -766 -535 -606
rect -496 -754 -490 -526
rect -456 -754 -450 -526
rect -398 -606 -392 -378
rect -358 -606 -352 -378
rect -313 -526 -303 -366
rect -251 -526 -241 -366
rect -202 -378 -156 -366
rect -496 -766 -450 -754
rect -411 -766 -401 -606
rect -349 -766 -339 -606
rect -300 -754 -294 -526
rect -260 -754 -254 -526
rect -202 -606 -196 -378
rect -162 -606 -156 -378
rect -117 -526 -107 -366
rect -55 -526 -45 -366
rect -6 -378 40 -366
rect -300 -766 -254 -754
rect -215 -766 -205 -606
rect -153 -766 -143 -606
rect -104 -754 -98 -526
rect -64 -754 -58 -526
rect -6 -606 0 -378
rect 34 -606 40 -378
rect 79 -526 89 -366
rect 141 -526 151 -366
rect 190 -378 236 -366
rect -104 -766 -58 -754
rect -19 -766 -9 -606
rect 43 -766 53 -606
rect 92 -754 98 -526
rect 132 -754 138 -526
rect 190 -606 196 -378
rect 230 -606 236 -378
rect 275 -526 285 -366
rect 337 -526 347 -366
rect 386 -378 432 -366
rect 92 -766 138 -754
rect 177 -766 187 -606
rect 239 -766 249 -606
rect 288 -754 294 -526
rect 328 -754 334 -526
rect 386 -606 392 -378
rect 426 -606 432 -378
rect 471 -526 481 -366
rect 533 -526 543 -366
rect 582 -378 628 -366
rect 288 -766 334 -754
rect 373 -766 383 -606
rect 435 -766 445 -606
rect 484 -754 490 -526
rect 524 -754 530 -526
rect 582 -606 588 -378
rect 622 -606 628 -378
rect 667 -526 677 -366
rect 729 -526 739 -366
rect 778 -378 824 -366
rect 484 -766 530 -754
rect 569 -766 579 -606
rect 631 -766 641 -606
rect 680 -754 686 -526
rect 720 -754 726 -526
rect 778 -606 784 -378
rect 818 -606 824 -378
rect 863 -526 873 -366
rect 925 -526 935 -366
rect 974 -378 1020 -366
rect 680 -766 726 -754
rect 765 -766 775 -606
rect 827 -766 837 -606
rect 876 -754 882 -526
rect 916 -754 922 -526
rect 974 -606 980 -378
rect 1014 -606 1020 -378
rect 1059 -526 1069 -366
rect 1121 -526 1131 -366
rect 1170 -378 1216 -366
rect 876 -766 922 -754
rect 961 -766 971 -606
rect 1023 -766 1033 -606
rect 1072 -754 1078 -526
rect 1112 -754 1118 -526
rect 1170 -606 1176 -378
rect 1210 -606 1216 -378
rect 1255 -526 1265 -366
rect 1317 -526 1327 -366
rect 1072 -766 1118 -754
rect 1157 -766 1167 -606
rect 1219 -766 1229 -606
rect 1268 -754 1274 -526
rect 1308 -754 1314 -526
rect 1268 -766 1314 -754
rect -1144 -800 1274 -794
rect 1404 -800 1544 -330
rect 2344 -290 2434 180
rect 2517 178 2533 180
rect 2567 178 2631 212
rect 2665 178 2729 212
rect 2763 178 2827 212
rect 2861 178 2925 212
rect 2959 178 3023 212
rect 3057 178 3121 212
rect 3155 178 3219 212
rect 3253 178 3317 212
rect 3351 178 3415 212
rect 3449 178 3513 212
rect 3547 178 3611 212
rect 3645 178 3709 212
rect 3743 178 3807 212
rect 3841 178 3905 212
rect 3939 178 3955 212
rect 2517 172 3955 178
rect 2478 128 2524 140
rect 2478 -100 2484 128
rect 2518 -100 2524 128
rect 2563 -20 2573 140
rect 2625 -20 2635 140
rect 2674 128 2720 140
rect 2465 -260 2475 -100
rect 2527 -260 2537 -100
rect 2576 -248 2582 -20
rect 2616 -248 2622 -20
rect 2674 -100 2680 128
rect 2714 -100 2720 128
rect 2759 -20 2769 140
rect 2821 -20 2831 140
rect 2870 128 2916 140
rect 2576 -260 2622 -248
rect 2661 -260 2671 -100
rect 2723 -260 2733 -100
rect 2772 -248 2778 -20
rect 2812 -248 2818 -20
rect 2870 -100 2876 128
rect 2910 -100 2916 128
rect 2955 -20 2965 140
rect 3017 -20 3027 140
rect 3066 128 3112 140
rect 2772 -260 2818 -248
rect 2857 -260 2867 -100
rect 2919 -260 2929 -100
rect 2968 -248 2974 -20
rect 3008 -248 3014 -20
rect 3066 -100 3072 128
rect 3106 -100 3112 128
rect 3151 -20 3161 140
rect 3213 -20 3223 140
rect 3262 128 3308 140
rect 2968 -260 3014 -248
rect 3053 -260 3063 -100
rect 3115 -260 3125 -100
rect 3164 -248 3170 -20
rect 3204 -248 3210 -20
rect 3262 -100 3268 128
rect 3302 -100 3308 128
rect 3347 -20 3357 140
rect 3409 -20 3419 140
rect 3458 128 3504 140
rect 3164 -260 3210 -248
rect 3249 -260 3259 -100
rect 3311 -260 3321 -100
rect 3360 -248 3366 -20
rect 3400 -248 3406 -20
rect 3458 -100 3464 128
rect 3498 -100 3504 128
rect 3543 -20 3553 140
rect 3605 -20 3615 140
rect 3654 128 3700 140
rect 3360 -260 3406 -248
rect 3445 -260 3455 -100
rect 3507 -260 3517 -100
rect 3556 -248 3562 -20
rect 3596 -248 3602 -20
rect 3654 -100 3660 128
rect 3694 -100 3700 128
rect 3739 -20 3749 140
rect 3801 -20 3811 140
rect 3850 128 3896 140
rect 3556 -260 3602 -248
rect 3641 -260 3651 -100
rect 3703 -260 3713 -100
rect 3752 -248 3758 -20
rect 3792 -248 3798 -20
rect 3850 -100 3856 128
rect 3890 -100 3896 128
rect 3935 -20 3945 140
rect 3997 -20 4007 140
rect 4044 130 4054 340
rect 4174 130 4184 340
rect 4048 118 4180 130
rect 3752 -260 3798 -248
rect 3837 -260 3847 -100
rect 3899 -260 3909 -100
rect 3948 -248 3954 -20
rect 3988 -248 3994 -20
rect 3948 -260 3994 -248
rect 2344 -292 2524 -290
rect 2344 -298 3955 -292
rect 2344 -332 2533 -298
rect 2567 -332 2631 -298
rect 2665 -332 2729 -298
rect 2763 -332 2827 -298
rect 2861 -332 2925 -298
rect 2959 -332 3023 -298
rect 3057 -332 3121 -298
rect 3155 -332 3219 -298
rect 3253 -332 3317 -298
rect 3351 -332 3415 -298
rect 3449 -332 3513 -298
rect 3547 -332 3611 -298
rect 3645 -332 3709 -298
rect 3743 -332 3807 -298
rect 3841 -332 3905 -298
rect 3939 -332 3955 -298
rect 2344 -348 3955 -332
rect 2344 -350 2524 -348
rect -1386 -804 1544 -800
rect -1386 -838 -1128 -804
rect -1094 -838 -1029 -804
rect -995 -838 -932 -804
rect -898 -838 -833 -804
rect -799 -838 -736 -804
rect -702 -838 -637 -804
rect -603 -838 -540 -804
rect -506 -838 -441 -804
rect -407 -838 -344 -804
rect -310 -838 -245 -804
rect -211 -838 -148 -804
rect -114 -838 -49 -804
rect -15 -838 48 -804
rect 82 -838 147 -804
rect 181 -838 244 -804
rect 278 -838 343 -804
rect 377 -838 440 -804
rect 474 -838 539 -804
rect 573 -838 636 -804
rect 670 -838 735 -804
rect 769 -838 832 -804
rect 866 -838 931 -804
rect 965 -838 1028 -804
rect 1062 -838 1127 -804
rect 1161 -838 1224 -804
rect 1258 -838 1544 -804
rect -1386 -912 1544 -838
rect -1386 -946 -1127 -912
rect -1093 -946 -1029 -912
rect -995 -946 -931 -912
rect -897 -946 -833 -912
rect -799 -946 -735 -912
rect -701 -946 -637 -912
rect -603 -946 -539 -912
rect -505 -946 -441 -912
rect -407 -946 -343 -912
rect -309 -946 -245 -912
rect -211 -946 -147 -912
rect -113 -946 -49 -912
rect -15 -946 49 -912
rect 83 -946 147 -912
rect 181 -946 245 -912
rect 279 -946 343 -912
rect 377 -946 441 -912
rect 475 -946 539 -912
rect 573 -946 637 -912
rect 671 -946 735 -912
rect 769 -946 833 -912
rect 867 -946 931 -912
rect 965 -946 1029 -912
rect 1063 -946 1127 -912
rect 1161 -946 1225 -912
rect 1259 -946 1544 -912
rect -1386 -950 1544 -946
rect -1386 -1020 -1236 -950
rect -1143 -956 1275 -950
rect -1860 -1260 -1236 -1020
rect -1195 -1144 -1185 -984
rect -1133 -1144 -1123 -984
rect -1084 -996 -1038 -984
rect -1386 -1420 -1236 -1260
rect -1182 -1372 -1176 -1144
rect -1142 -1372 -1136 -1144
rect -1084 -1224 -1078 -996
rect -1044 -1224 -1038 -996
rect -999 -1144 -989 -984
rect -937 -1144 -927 -984
rect -888 -996 -842 -984
rect -1182 -1384 -1136 -1372
rect -1097 -1384 -1087 -1224
rect -1035 -1384 -1025 -1224
rect -986 -1372 -980 -1144
rect -946 -1372 -940 -1144
rect -888 -1224 -882 -996
rect -848 -1224 -842 -996
rect -803 -1144 -793 -984
rect -741 -1144 -731 -984
rect -692 -996 -646 -984
rect -986 -1384 -940 -1372
rect -901 -1384 -891 -1224
rect -839 -1384 -829 -1224
rect -790 -1372 -784 -1144
rect -750 -1372 -744 -1144
rect -692 -1224 -686 -996
rect -652 -1224 -646 -996
rect -607 -1144 -597 -984
rect -545 -1144 -535 -984
rect -496 -996 -450 -984
rect -790 -1384 -744 -1372
rect -705 -1384 -695 -1224
rect -643 -1384 -633 -1224
rect -594 -1372 -588 -1144
rect -554 -1372 -548 -1144
rect -496 -1224 -490 -996
rect -456 -1224 -450 -996
rect -411 -1144 -401 -984
rect -349 -1144 -339 -984
rect -300 -996 -254 -984
rect -594 -1384 -548 -1372
rect -509 -1384 -499 -1224
rect -447 -1384 -437 -1224
rect -398 -1372 -392 -1144
rect -358 -1372 -352 -1144
rect -300 -1224 -294 -996
rect -260 -1224 -254 -996
rect -215 -1144 -205 -984
rect -153 -1144 -143 -984
rect -104 -996 -58 -984
rect -398 -1384 -352 -1372
rect -313 -1384 -303 -1224
rect -251 -1384 -241 -1224
rect -202 -1372 -196 -1144
rect -162 -1372 -156 -1144
rect -104 -1224 -98 -996
rect -64 -1224 -58 -996
rect -19 -1144 -9 -984
rect 43 -1144 53 -984
rect 92 -996 138 -984
rect -202 -1384 -156 -1372
rect -117 -1384 -107 -1224
rect -55 -1384 -45 -1224
rect -6 -1372 0 -1144
rect 34 -1372 40 -1144
rect 92 -1224 98 -996
rect 132 -1224 138 -996
rect 177 -1144 187 -984
rect 239 -1144 249 -984
rect 288 -996 334 -984
rect -6 -1384 40 -1372
rect 79 -1384 89 -1224
rect 141 -1384 151 -1224
rect 190 -1372 196 -1144
rect 230 -1372 236 -1144
rect 288 -1224 294 -996
rect 328 -1224 334 -996
rect 373 -1144 383 -984
rect 435 -1144 445 -984
rect 484 -996 530 -984
rect 190 -1384 236 -1372
rect 275 -1384 285 -1224
rect 337 -1384 347 -1224
rect 386 -1372 392 -1144
rect 426 -1372 432 -1144
rect 484 -1224 490 -996
rect 524 -1224 530 -996
rect 569 -1144 579 -984
rect 631 -1144 641 -984
rect 680 -996 726 -984
rect 386 -1384 432 -1372
rect 471 -1384 481 -1224
rect 533 -1384 543 -1224
rect 582 -1372 588 -1144
rect 622 -1372 628 -1144
rect 680 -1224 686 -996
rect 720 -1224 726 -996
rect 765 -1144 775 -984
rect 827 -1144 837 -984
rect 876 -996 922 -984
rect 582 -1384 628 -1372
rect 667 -1384 677 -1224
rect 729 -1384 739 -1224
rect 778 -1372 784 -1144
rect 818 -1372 824 -1144
rect 876 -1224 882 -996
rect 916 -1224 922 -996
rect 961 -1144 971 -984
rect 1023 -1144 1033 -984
rect 1072 -996 1118 -984
rect 778 -1384 824 -1372
rect 863 -1384 873 -1224
rect 925 -1384 935 -1224
rect 974 -1372 980 -1144
rect 1014 -1372 1020 -1144
rect 1072 -1224 1078 -996
rect 1112 -1224 1118 -996
rect 1157 -1144 1167 -984
rect 1219 -1144 1229 -984
rect 1268 -996 1314 -984
rect 974 -1384 1020 -1372
rect 1059 -1384 1069 -1224
rect 1121 -1384 1131 -1224
rect 1170 -1372 1176 -1144
rect 1210 -1372 1216 -1144
rect 1268 -1224 1274 -996
rect 1308 -1224 1314 -996
rect 1170 -1384 1216 -1372
rect 1255 -1384 1265 -1224
rect 1317 -1384 1327 -1224
rect 1404 -1410 1544 -950
rect 1644 -948 2964 -920
rect 1644 -982 1662 -948
rect 1696 -982 1758 -948
rect 1792 -982 1854 -948
rect 1888 -982 1950 -948
rect 1984 -982 2046 -948
rect 2080 -982 2142 -948
rect 2176 -982 2238 -948
rect 2272 -982 2334 -948
rect 2368 -982 2430 -948
rect 2464 -982 2526 -948
rect 2560 -982 2622 -948
rect 2656 -982 2718 -948
rect 2752 -982 2964 -948
rect 1644 -990 2964 -982
rect 1608 -1032 1654 -1020
rect 1608 -1260 1614 -1032
rect 1648 -1260 1654 -1032
rect 1691 -1180 1701 -1020
rect 1753 -1180 1763 -1020
rect 1800 -1032 1846 -1020
rect -1143 -1420 1275 -1412
rect 1384 -1420 1544 -1410
rect 1595 -1420 1605 -1260
rect 1657 -1420 1667 -1260
rect 1704 -1408 1710 -1180
rect 1744 -1408 1750 -1180
rect 1800 -1260 1806 -1032
rect 1840 -1260 1846 -1032
rect 1883 -1180 1893 -1020
rect 1945 -1180 1955 -1020
rect 1992 -1032 2038 -1020
rect 1704 -1420 1750 -1408
rect 1787 -1420 1797 -1260
rect 1849 -1420 1859 -1260
rect 1896 -1408 1902 -1180
rect 1936 -1408 1942 -1180
rect 1992 -1260 1998 -1032
rect 2032 -1260 2038 -1032
rect 2075 -1180 2085 -1020
rect 2137 -1180 2147 -1020
rect 2184 -1032 2230 -1020
rect 1896 -1420 1942 -1408
rect 1979 -1420 1989 -1260
rect 2041 -1420 2051 -1260
rect 2088 -1408 2094 -1180
rect 2128 -1408 2134 -1180
rect 2184 -1260 2190 -1032
rect 2224 -1260 2230 -1032
rect 2267 -1180 2277 -1020
rect 2329 -1180 2339 -1020
rect 2376 -1032 2422 -1020
rect 2088 -1420 2134 -1408
rect 2171 -1420 2181 -1260
rect 2233 -1420 2243 -1260
rect 2280 -1408 2286 -1180
rect 2320 -1408 2326 -1180
rect 2376 -1260 2382 -1032
rect 2416 -1260 2422 -1032
rect 2459 -1180 2469 -1020
rect 2521 -1180 2531 -1020
rect 2568 -1032 2614 -1020
rect 2280 -1420 2326 -1408
rect 2363 -1420 2373 -1260
rect 2425 -1420 2435 -1260
rect 2472 -1408 2478 -1180
rect 2512 -1408 2518 -1180
rect 2568 -1260 2574 -1032
rect 2608 -1260 2614 -1032
rect 2651 -1180 2661 -1020
rect 2713 -1180 2723 -1020
rect 2760 -1032 2806 -1020
rect 2472 -1420 2518 -1408
rect 2555 -1420 2565 -1260
rect 2617 -1420 2627 -1260
rect 2664 -1408 2670 -1180
rect 2704 -1408 2710 -1180
rect 2760 -1260 2766 -1032
rect 2800 -1260 2806 -1032
rect 2664 -1420 2710 -1408
rect 2747 -1420 2757 -1260
rect 2809 -1420 2819 -1260
rect -1386 -1422 1544 -1420
rect -1386 -1456 -1127 -1422
rect -1093 -1456 -1029 -1422
rect -995 -1456 -931 -1422
rect -897 -1456 -833 -1422
rect -799 -1456 -735 -1422
rect -701 -1456 -637 -1422
rect -603 -1456 -539 -1422
rect -505 -1456 -441 -1422
rect -407 -1456 -343 -1422
rect -309 -1456 -245 -1422
rect -211 -1456 -147 -1422
rect -113 -1456 -49 -1422
rect -15 -1456 49 -1422
rect 83 -1456 147 -1422
rect 181 -1456 245 -1422
rect 279 -1456 343 -1422
rect 377 -1456 441 -1422
rect 475 -1456 539 -1422
rect 573 -1456 637 -1422
rect 671 -1456 735 -1422
rect 769 -1456 833 -1422
rect 867 -1456 931 -1422
rect 965 -1456 1029 -1422
rect 1063 -1456 1127 -1422
rect 1161 -1456 1225 -1422
rect 1259 -1456 1544 -1422
rect 2854 -1450 2964 -990
rect -1386 -1470 1544 -1456
rect 1644 -1458 2964 -1450
rect -1143 -1472 1275 -1470
rect 1644 -1492 1662 -1458
rect 1696 -1492 1758 -1458
rect 1792 -1492 1854 -1458
rect 1888 -1492 1950 -1458
rect 1984 -1492 2046 -1458
rect 2080 -1492 2142 -1458
rect 2176 -1492 2238 -1458
rect 2272 -1492 2334 -1458
rect 2368 -1492 2430 -1458
rect 2464 -1492 2526 -1458
rect 2560 -1492 2622 -1458
rect 2656 -1492 2718 -1458
rect 2752 -1492 2964 -1458
rect 1644 -1520 2964 -1492
rect 2834 -1660 2964 -1520
rect -1346 -1697 -1196 -1690
rect -1346 -1714 1247 -1697
rect -1346 -1748 -1148 -1714
rect -1114 -1748 -956 -1714
rect -922 -1748 -764 -1714
rect -730 -1748 -572 -1714
rect -538 -1748 -380 -1714
rect -346 -1748 -188 -1714
rect -154 -1748 4 -1714
rect 38 -1748 196 -1714
rect 230 -1748 388 -1714
rect 422 -1748 580 -1714
rect 614 -1748 772 -1714
rect 806 -1748 964 -1714
rect 998 -1748 1156 -1714
rect 1190 -1748 1247 -1714
rect 2834 -1730 3140 -1660
rect -1346 -1750 1247 -1748
rect -1346 -2220 -1246 -1750
rect -1203 -1757 1247 -1750
rect 1654 -1768 3140 -1730
rect -1202 -1798 -1156 -1786
rect -1202 -2026 -1196 -1798
rect -1162 -2026 -1156 -1798
rect -1119 -1946 -1109 -1786
rect -1057 -1946 -1047 -1786
rect -1010 -1798 -964 -1786
rect -1215 -2186 -1205 -2026
rect -1153 -2186 -1143 -2026
rect -1106 -2174 -1100 -1946
rect -1066 -2174 -1060 -1946
rect -1010 -2026 -1004 -1798
rect -970 -2026 -964 -1798
rect -927 -1946 -917 -1786
rect -865 -1946 -855 -1786
rect -818 -1798 -772 -1786
rect -1106 -2186 -1060 -2174
rect -1023 -2186 -1013 -2026
rect -961 -2186 -951 -2026
rect -914 -2174 -908 -1946
rect -874 -2174 -868 -1946
rect -818 -2026 -812 -1798
rect -778 -2026 -772 -1798
rect -735 -1946 -725 -1786
rect -673 -1946 -663 -1786
rect -626 -1798 -580 -1786
rect -914 -2186 -868 -2174
rect -831 -2186 -821 -2026
rect -769 -2186 -759 -2026
rect -722 -2174 -716 -1946
rect -682 -2174 -676 -1946
rect -626 -2026 -620 -1798
rect -586 -2026 -580 -1798
rect -543 -1946 -533 -1786
rect -481 -1946 -471 -1786
rect -434 -1798 -388 -1786
rect -722 -2186 -676 -2174
rect -639 -2186 -629 -2026
rect -577 -2186 -567 -2026
rect -530 -2174 -524 -1946
rect -490 -2174 -484 -1946
rect -434 -2026 -428 -1798
rect -394 -2026 -388 -1798
rect -351 -1946 -341 -1786
rect -289 -1946 -279 -1786
rect -242 -1798 -196 -1786
rect -530 -2186 -484 -2174
rect -447 -2186 -437 -2026
rect -385 -2186 -375 -2026
rect -338 -2174 -332 -1946
rect -298 -2174 -292 -1946
rect -242 -2026 -236 -1798
rect -202 -2026 -196 -1798
rect -159 -1946 -149 -1786
rect -97 -1946 -87 -1786
rect -50 -1798 -4 -1786
rect -338 -2186 -292 -2174
rect -255 -2186 -245 -2026
rect -193 -2186 -183 -2026
rect -146 -2174 -140 -1946
rect -106 -2174 -100 -1946
rect -50 -2026 -44 -1798
rect -10 -2026 -4 -1798
rect 33 -1946 43 -1786
rect 95 -1946 105 -1786
rect 142 -1798 188 -1786
rect -146 -2186 -100 -2174
rect -63 -2186 -53 -2026
rect -1 -2186 9 -2026
rect 46 -2174 52 -1946
rect 86 -2174 92 -1946
rect 142 -2026 148 -1798
rect 182 -2026 188 -1798
rect 225 -1946 235 -1786
rect 287 -1946 297 -1786
rect 334 -1798 380 -1786
rect 46 -2186 92 -2174
rect 129 -2186 139 -2026
rect 191 -2186 201 -2026
rect 238 -2174 244 -1946
rect 278 -2174 284 -1946
rect 334 -2026 340 -1798
rect 374 -2026 380 -1798
rect 417 -1946 427 -1786
rect 479 -1946 489 -1786
rect 526 -1798 572 -1786
rect 238 -2186 284 -2174
rect 321 -2186 331 -2026
rect 383 -2186 393 -2026
rect 430 -2174 436 -1946
rect 470 -2174 476 -1946
rect 526 -2026 532 -1798
rect 566 -2026 572 -1798
rect 609 -1946 619 -1786
rect 671 -1946 681 -1786
rect 718 -1798 764 -1786
rect 430 -2186 476 -2174
rect 513 -2186 523 -2026
rect 575 -2186 585 -2026
rect 622 -2174 628 -1946
rect 662 -2174 668 -1946
rect 718 -2026 724 -1798
rect 758 -2026 764 -1798
rect 801 -1946 811 -1786
rect 863 -1946 873 -1786
rect 910 -1798 956 -1786
rect 622 -2186 668 -2174
rect 705 -2186 715 -2026
rect 767 -2186 777 -2026
rect 814 -2174 820 -1946
rect 854 -2174 860 -1946
rect 910 -2026 916 -1798
rect 950 -2026 956 -1798
rect 993 -1946 1003 -1786
rect 1055 -1946 1065 -1786
rect 1102 -1798 1148 -1786
rect 814 -2186 860 -2174
rect 897 -2186 907 -2026
rect 959 -2186 969 -2026
rect 1006 -2174 1012 -1946
rect 1046 -2174 1052 -1946
rect 1102 -2026 1108 -1798
rect 1142 -2026 1148 -1798
rect 1185 -1946 1195 -1786
rect 1247 -1946 1257 -1786
rect 1654 -1802 1676 -1768
rect 1844 -1802 1934 -1768
rect 2102 -1802 2192 -1768
rect 2360 -1802 2450 -1768
rect 2618 -1802 2708 -1768
rect 2876 -1802 2966 -1768
rect 3134 -1780 3140 -1768
rect 3320 -1780 3330 -1660
rect 3134 -1802 3330 -1780
rect 1654 -1810 3330 -1802
rect 1608 -1852 1654 -1840
rect 1006 -2186 1052 -2174
rect 1089 -2186 1099 -2026
rect 1151 -2186 1161 -2026
rect 1198 -2174 1204 -1946
rect 1238 -2174 1244 -1946
rect 1338 -2070 1480 -2058
rect 1198 -2186 1244 -2174
rect -1203 -2220 1247 -2217
rect -1346 -2224 1247 -2220
rect -1346 -2258 -1052 -2224
rect -1018 -2258 -860 -2224
rect -826 -2258 -668 -2224
rect -634 -2258 -476 -2224
rect -442 -2258 -284 -2224
rect -250 -2258 -92 -2224
rect -58 -2258 100 -2224
rect 134 -2258 292 -2224
rect 326 -2258 484 -2224
rect 518 -2258 676 -2224
rect 710 -2258 868 -2224
rect 902 -2258 1060 -2224
rect 1094 -2258 1247 -2224
rect 1334 -2250 1344 -2070
rect 1474 -2250 1484 -2070
rect 1608 -2080 1614 -1852
rect 1648 -2080 1654 -1852
rect 1853 -2000 1863 -1840
rect 1915 -2000 1925 -1840
rect 2124 -1852 2170 -1840
rect 1595 -2240 1605 -2080
rect 1657 -2240 1667 -2080
rect 1866 -2228 1872 -2000
rect 1906 -2228 1912 -2000
rect 2124 -2080 2130 -1852
rect 2164 -2080 2170 -1852
rect 2369 -2000 2379 -1840
rect 2431 -2000 2441 -1840
rect 2640 -1852 2686 -1840
rect 1866 -2240 1912 -2228
rect 2111 -2240 2121 -2080
rect 2173 -2240 2183 -2080
rect 2382 -2228 2388 -2000
rect 2422 -2228 2428 -2000
rect 2640 -2080 2646 -1852
rect 2680 -2080 2686 -1852
rect 2885 -2000 2895 -1840
rect 2947 -2000 2954 -1840
rect 2382 -2240 2428 -2228
rect 2627 -2240 2637 -2080
rect 2689 -2240 2699 -2080
rect 2898 -2228 2904 -2000
rect 2938 -2228 2944 -2000
rect 2898 -2240 2944 -2228
rect -1346 -2332 1247 -2258
rect 1338 -2262 1480 -2250
rect 3004 -2270 3094 -1810
rect 3156 -1852 3202 -1840
rect 3156 -2080 3162 -1852
rect 3196 -2080 3202 -1852
rect 3143 -2240 3153 -2080
rect 3205 -2240 3215 -2080
rect -1346 -2366 -1052 -2332
rect -1018 -2366 -860 -2332
rect -826 -2366 -668 -2332
rect -634 -2366 -476 -2332
rect -442 -2366 -284 -2332
rect -250 -2366 -92 -2332
rect -58 -2366 100 -2332
rect 134 -2366 292 -2332
rect 326 -2366 484 -2332
rect 518 -2366 676 -2332
rect 710 -2366 868 -2332
rect 902 -2366 1060 -2332
rect 1094 -2366 1247 -2332
rect 1594 -2278 4620 -2270
rect 1594 -2312 1676 -2278
rect 1844 -2312 1934 -2278
rect 2102 -2312 2192 -2278
rect 2360 -2312 2450 -2278
rect 2618 -2312 2708 -2278
rect 2876 -2312 2966 -2278
rect 3134 -2312 4620 -2278
rect 1594 -2350 4620 -2312
rect -1346 -2367 1247 -2366
rect -1346 -2370 -1196 -2367
rect -1346 -2840 -1246 -2370
rect -1064 -2372 -1006 -2367
rect -872 -2372 -814 -2367
rect -680 -2372 -622 -2367
rect -488 -2372 -430 -2367
rect -296 -2372 -238 -2367
rect -104 -2372 -46 -2367
rect 88 -2372 146 -2367
rect 280 -2372 338 -2367
rect 472 -2372 530 -2367
rect 664 -2372 722 -2367
rect 856 -2372 914 -2367
rect 1048 -2372 1106 -2367
rect -1215 -2564 -1205 -2404
rect -1153 -2564 -1143 -2404
rect -1106 -2416 -1060 -2404
rect -1202 -2792 -1196 -2564
rect -1162 -2792 -1156 -2564
rect -1106 -2644 -1100 -2416
rect -1066 -2644 -1060 -2416
rect -1023 -2564 -1013 -2404
rect -961 -2564 -951 -2404
rect -914 -2416 -868 -2404
rect -1202 -2804 -1156 -2792
rect -1119 -2804 -1109 -2644
rect -1057 -2804 -1047 -2644
rect -1010 -2792 -1004 -2564
rect -970 -2792 -964 -2564
rect -914 -2644 -908 -2416
rect -874 -2644 -868 -2416
rect -831 -2564 -821 -2404
rect -769 -2564 -759 -2404
rect -722 -2416 -676 -2404
rect -1010 -2804 -964 -2792
rect -927 -2804 -917 -2644
rect -865 -2804 -855 -2644
rect -818 -2792 -812 -2564
rect -778 -2792 -772 -2564
rect -722 -2644 -716 -2416
rect -682 -2644 -676 -2416
rect -639 -2564 -629 -2404
rect -577 -2564 -567 -2404
rect -530 -2416 -484 -2404
rect -818 -2804 -772 -2792
rect -735 -2804 -725 -2644
rect -673 -2804 -663 -2644
rect -626 -2792 -620 -2564
rect -586 -2792 -580 -2564
rect -530 -2644 -524 -2416
rect -490 -2644 -484 -2416
rect -447 -2564 -437 -2404
rect -385 -2564 -375 -2404
rect -338 -2416 -292 -2404
rect -626 -2804 -580 -2792
rect -543 -2804 -533 -2644
rect -481 -2804 -471 -2644
rect -434 -2792 -428 -2564
rect -394 -2792 -388 -2564
rect -338 -2644 -332 -2416
rect -298 -2644 -292 -2416
rect -255 -2564 -245 -2404
rect -193 -2564 -183 -2404
rect -146 -2416 -100 -2404
rect -434 -2804 -388 -2792
rect -351 -2804 -341 -2644
rect -289 -2804 -279 -2644
rect -242 -2792 -236 -2564
rect -202 -2792 -196 -2564
rect -146 -2644 -140 -2416
rect -106 -2644 -100 -2416
rect -63 -2564 -53 -2404
rect -1 -2564 9 -2404
rect 46 -2416 92 -2404
rect -242 -2804 -196 -2792
rect -159 -2804 -149 -2644
rect -97 -2804 -87 -2644
rect -50 -2792 -44 -2564
rect -10 -2792 -4 -2564
rect 46 -2644 52 -2416
rect 86 -2644 92 -2416
rect 129 -2564 139 -2404
rect 191 -2564 201 -2404
rect 238 -2416 284 -2404
rect -50 -2804 -4 -2792
rect 33 -2804 43 -2644
rect 95 -2804 105 -2644
rect 142 -2792 148 -2564
rect 182 -2792 188 -2564
rect 238 -2644 244 -2416
rect 278 -2644 284 -2416
rect 321 -2564 331 -2404
rect 383 -2564 393 -2404
rect 430 -2416 476 -2404
rect 142 -2804 188 -2792
rect 225 -2804 235 -2644
rect 287 -2804 297 -2644
rect 334 -2792 340 -2564
rect 374 -2792 380 -2564
rect 430 -2644 436 -2416
rect 470 -2644 476 -2416
rect 513 -2564 523 -2404
rect 575 -2564 585 -2404
rect 622 -2416 668 -2404
rect 334 -2804 380 -2792
rect 417 -2804 427 -2644
rect 479 -2804 489 -2644
rect 526 -2792 532 -2564
rect 566 -2792 572 -2564
rect 622 -2644 628 -2416
rect 662 -2644 668 -2416
rect 705 -2564 715 -2404
rect 767 -2564 777 -2404
rect 814 -2416 860 -2404
rect 526 -2804 572 -2792
rect 609 -2804 619 -2644
rect 671 -2804 681 -2644
rect 718 -2792 724 -2564
rect 758 -2792 764 -2564
rect 814 -2644 820 -2416
rect 854 -2644 860 -2416
rect 897 -2564 907 -2404
rect 959 -2564 969 -2404
rect 1006 -2416 1052 -2404
rect 718 -2804 764 -2792
rect 801 -2804 811 -2644
rect 863 -2804 873 -2644
rect 910 -2792 916 -2564
rect 950 -2792 956 -2564
rect 1006 -2644 1012 -2416
rect 1046 -2644 1052 -2416
rect 1089 -2564 1099 -2404
rect 1151 -2564 1161 -2404
rect 1198 -2416 1244 -2404
rect 910 -2804 956 -2792
rect 993 -2804 1003 -2644
rect 1055 -2804 1065 -2644
rect 1102 -2792 1108 -2564
rect 1142 -2792 1148 -2564
rect 1198 -2644 1204 -2416
rect 1238 -2644 1244 -2416
rect 1102 -2804 1148 -2792
rect 1185 -2804 1195 -2644
rect 1247 -2804 1257 -2644
rect -1160 -2837 -1102 -2836
rect -968 -2837 -910 -2836
rect -776 -2837 -718 -2836
rect -584 -2837 -526 -2836
rect -392 -2837 -334 -2836
rect -200 -2837 -142 -2836
rect -8 -2837 50 -2836
rect 184 -2837 242 -2836
rect 376 -2837 434 -2836
rect 568 -2837 626 -2836
rect 760 -2837 818 -2836
rect 952 -2837 1010 -2836
rect 1144 -2837 1202 -2836
rect -1203 -2840 1247 -2837
rect -1346 -2842 1247 -2840
rect -1346 -2876 -1148 -2842
rect -1114 -2876 -956 -2842
rect -922 -2876 -764 -2842
rect -730 -2876 -572 -2842
rect -538 -2876 -380 -2842
rect -346 -2876 -188 -2842
rect -154 -2876 4 -2842
rect 38 -2876 196 -2842
rect 230 -2876 388 -2842
rect 422 -2876 580 -2842
rect 614 -2876 772 -2842
rect 806 -2876 964 -2842
rect 998 -2876 1156 -2842
rect 1190 -2876 1247 -2842
rect -1346 -2950 1247 -2876
rect -1346 -2984 -1148 -2950
rect -1114 -2984 -956 -2950
rect -922 -2984 -764 -2950
rect -730 -2984 -572 -2950
rect -538 -2984 -380 -2950
rect -346 -2984 -188 -2950
rect -154 -2984 4 -2950
rect 38 -2984 196 -2950
rect 230 -2984 388 -2950
rect 422 -2984 580 -2950
rect 614 -2984 772 -2950
rect 806 -2984 964 -2950
rect 998 -2984 1156 -2950
rect 1190 -2984 1247 -2950
rect -1346 -2987 1247 -2984
rect -1346 -2990 -1102 -2987
rect -968 -2990 -910 -2987
rect -776 -2990 -718 -2987
rect -584 -2990 -526 -2987
rect -392 -2990 -334 -2987
rect -200 -2990 -142 -2987
rect -8 -2990 50 -2987
rect 184 -2990 242 -2987
rect 376 -2990 434 -2987
rect 568 -2990 626 -2987
rect 760 -2990 818 -2987
rect 952 -2990 1010 -2987
rect 1144 -2990 1202 -2987
rect -1346 -3460 -1246 -2990
rect -1202 -3034 -1156 -3022
rect -1202 -3262 -1196 -3034
rect -1162 -3262 -1156 -3034
rect -1119 -3182 -1109 -3022
rect -1057 -3182 -1047 -3022
rect -1010 -3034 -964 -3022
rect -1215 -3422 -1205 -3262
rect -1153 -3422 -1143 -3262
rect -1106 -3410 -1100 -3182
rect -1066 -3410 -1060 -3182
rect -1010 -3262 -1004 -3034
rect -970 -3262 -964 -3034
rect -927 -3182 -917 -3022
rect -865 -3182 -855 -3022
rect -818 -3034 -772 -3022
rect -1106 -3422 -1060 -3410
rect -1023 -3422 -1013 -3262
rect -961 -3422 -951 -3262
rect -914 -3410 -908 -3182
rect -874 -3410 -868 -3182
rect -818 -3262 -812 -3034
rect -778 -3262 -772 -3034
rect -735 -3182 -725 -3022
rect -673 -3182 -663 -3022
rect -626 -3034 -580 -3022
rect -914 -3422 -868 -3410
rect -831 -3422 -821 -3262
rect -769 -3422 -759 -3262
rect -722 -3410 -716 -3182
rect -682 -3410 -676 -3182
rect -626 -3262 -620 -3034
rect -586 -3262 -580 -3034
rect -543 -3182 -533 -3022
rect -481 -3182 -471 -3022
rect -434 -3034 -388 -3022
rect -722 -3422 -676 -3410
rect -639 -3422 -629 -3262
rect -577 -3422 -567 -3262
rect -530 -3410 -524 -3182
rect -490 -3410 -484 -3182
rect -434 -3262 -428 -3034
rect -394 -3262 -388 -3034
rect -351 -3182 -341 -3022
rect -289 -3182 -279 -3022
rect -242 -3034 -196 -3022
rect -530 -3422 -484 -3410
rect -447 -3422 -437 -3262
rect -385 -3422 -375 -3262
rect -338 -3410 -332 -3182
rect -298 -3410 -292 -3182
rect -242 -3262 -236 -3034
rect -202 -3262 -196 -3034
rect -159 -3182 -149 -3022
rect -97 -3182 -87 -3022
rect -50 -3034 -4 -3022
rect -338 -3422 -292 -3410
rect -255 -3422 -245 -3262
rect -193 -3422 -183 -3262
rect -146 -3410 -140 -3182
rect -106 -3410 -100 -3182
rect -50 -3262 -44 -3034
rect -10 -3262 -4 -3034
rect 33 -3182 43 -3022
rect 95 -3182 105 -3022
rect 142 -3034 188 -3022
rect -146 -3422 -100 -3410
rect -63 -3422 -53 -3262
rect -1 -3422 9 -3262
rect 46 -3410 52 -3182
rect 86 -3410 92 -3182
rect 142 -3262 148 -3034
rect 182 -3262 188 -3034
rect 225 -3182 235 -3022
rect 287 -3182 297 -3022
rect 334 -3034 380 -3022
rect 46 -3422 92 -3410
rect 129 -3422 139 -3262
rect 191 -3422 201 -3262
rect 238 -3410 244 -3182
rect 278 -3410 284 -3182
rect 334 -3262 340 -3034
rect 374 -3262 380 -3034
rect 417 -3182 427 -3022
rect 479 -3182 489 -3022
rect 526 -3034 572 -3022
rect 238 -3422 284 -3410
rect 321 -3422 331 -3262
rect 383 -3422 393 -3262
rect 430 -3410 436 -3182
rect 470 -3410 476 -3182
rect 526 -3262 532 -3034
rect 566 -3262 572 -3034
rect 609 -3182 619 -3022
rect 671 -3182 681 -3022
rect 718 -3034 764 -3022
rect 430 -3422 476 -3410
rect 513 -3422 523 -3262
rect 575 -3422 585 -3262
rect 622 -3410 628 -3182
rect 662 -3410 668 -3182
rect 718 -3262 724 -3034
rect 758 -3262 764 -3034
rect 801 -3182 811 -3022
rect 863 -3182 873 -3022
rect 910 -3034 956 -3022
rect 622 -3422 668 -3410
rect 705 -3422 715 -3262
rect 767 -3422 777 -3262
rect 814 -3410 820 -3182
rect 854 -3410 860 -3182
rect 910 -3262 916 -3034
rect 950 -3262 956 -3034
rect 993 -3182 1003 -3022
rect 1055 -3182 1065 -3022
rect 1102 -3034 1148 -3022
rect 814 -3422 860 -3410
rect 897 -3422 907 -3262
rect 959 -3422 969 -3262
rect 1006 -3410 1012 -3182
rect 1046 -3410 1052 -3182
rect 1102 -3262 1108 -3034
rect 1142 -3262 1148 -3034
rect 1185 -3182 1195 -3022
rect 1247 -3182 1257 -3022
rect 1006 -3422 1052 -3410
rect 1089 -3422 1099 -3262
rect 1151 -3422 1161 -3262
rect 1198 -3410 1204 -3182
rect 1238 -3410 1244 -3182
rect 1198 -3422 1244 -3410
rect -1064 -3457 -1006 -3454
rect -872 -3457 -814 -3454
rect -680 -3457 -622 -3454
rect -488 -3457 -430 -3454
rect -296 -3457 -238 -3454
rect -104 -3457 -46 -3454
rect 88 -3457 146 -3454
rect 280 -3457 338 -3454
rect 472 -3457 530 -3454
rect 664 -3457 722 -3454
rect 856 -3457 914 -3454
rect 1048 -3457 1106 -3454
rect -1203 -3460 1247 -3457
rect -1346 -3494 -1052 -3460
rect -1018 -3494 -860 -3460
rect -826 -3494 -668 -3460
rect -634 -3494 -476 -3460
rect -442 -3494 -284 -3460
rect -250 -3494 -92 -3460
rect -58 -3494 100 -3460
rect 134 -3494 292 -3460
rect 326 -3494 484 -3460
rect 518 -3494 676 -3460
rect 710 -3494 868 -3460
rect 902 -3494 1060 -3460
rect 1094 -3494 1247 -3460
rect -1346 -3568 1247 -3494
rect -1346 -3602 -1052 -3568
rect -1018 -3602 -860 -3568
rect -826 -3602 -668 -3568
rect -634 -3602 -476 -3568
rect -442 -3602 -284 -3568
rect -250 -3602 -92 -3568
rect -58 -3602 100 -3568
rect 134 -3602 292 -3568
rect 326 -3602 484 -3568
rect 518 -3602 676 -3568
rect 710 -3602 868 -3568
rect 902 -3602 1060 -3568
rect 1094 -3602 1247 -3568
rect -1346 -3607 1247 -3602
rect -1346 -3610 -1186 -3607
rect -1064 -3608 -1006 -3607
rect -872 -3608 -814 -3607
rect -680 -3608 -622 -3607
rect -488 -3608 -430 -3607
rect -296 -3608 -238 -3607
rect -104 -3608 -46 -3607
rect 88 -3608 146 -3607
rect 280 -3608 338 -3607
rect 472 -3608 530 -3607
rect 664 -3608 722 -3607
rect 856 -3608 914 -3607
rect 1048 -3608 1106 -3607
rect -1346 -4020 -1246 -3610
rect -1215 -3800 -1205 -3640
rect -1153 -3800 -1143 -3640
rect -1106 -3652 -1060 -3640
rect -1390 -4120 -1380 -4020
rect -1270 -4080 -1246 -4020
rect -1202 -4028 -1196 -3800
rect -1162 -4028 -1156 -3800
rect -1106 -3880 -1100 -3652
rect -1066 -3880 -1060 -3652
rect -1023 -3800 -1013 -3640
rect -961 -3800 -951 -3640
rect -914 -3652 -868 -3640
rect -1202 -4040 -1156 -4028
rect -1119 -4040 -1109 -3880
rect -1057 -4040 -1047 -3880
rect -1010 -4028 -1004 -3800
rect -970 -4028 -964 -3800
rect -914 -3880 -908 -3652
rect -874 -3880 -868 -3652
rect -831 -3800 -821 -3640
rect -769 -3800 -759 -3640
rect -722 -3652 -676 -3640
rect -1010 -4040 -964 -4028
rect -927 -4040 -917 -3880
rect -865 -4040 -855 -3880
rect -818 -4028 -812 -3800
rect -778 -4028 -772 -3800
rect -722 -3880 -716 -3652
rect -682 -3880 -676 -3652
rect -639 -3800 -629 -3640
rect -577 -3800 -567 -3640
rect -530 -3652 -484 -3640
rect -818 -4040 -772 -4028
rect -735 -4040 -725 -3880
rect -673 -4040 -663 -3880
rect -626 -4028 -620 -3800
rect -586 -4028 -580 -3800
rect -530 -3880 -524 -3652
rect -490 -3880 -484 -3652
rect -447 -3800 -437 -3640
rect -385 -3800 -375 -3640
rect -338 -3652 -292 -3640
rect -626 -4040 -580 -4028
rect -543 -4040 -533 -3880
rect -481 -4040 -471 -3880
rect -434 -4028 -428 -3800
rect -394 -4028 -388 -3800
rect -338 -3880 -332 -3652
rect -298 -3880 -292 -3652
rect -255 -3800 -245 -3640
rect -193 -3800 -183 -3640
rect -146 -3652 -100 -3640
rect -434 -4040 -388 -4028
rect -351 -4040 -341 -3880
rect -289 -4040 -279 -3880
rect -242 -4028 -236 -3800
rect -202 -4028 -196 -3800
rect -146 -3880 -140 -3652
rect -106 -3880 -100 -3652
rect -63 -3800 -53 -3640
rect -1 -3800 9 -3640
rect 46 -3652 92 -3640
rect -242 -4040 -196 -4028
rect -159 -4040 -149 -3880
rect -97 -4040 -87 -3880
rect -50 -4028 -44 -3800
rect -10 -4028 -4 -3800
rect 46 -3880 52 -3652
rect 86 -3880 92 -3652
rect 129 -3800 139 -3640
rect 191 -3800 201 -3640
rect 238 -3652 284 -3640
rect -50 -4040 -4 -4028
rect 33 -4040 43 -3880
rect 95 -4040 105 -3880
rect 142 -4028 148 -3800
rect 182 -4028 188 -3800
rect 238 -3880 244 -3652
rect 278 -3880 284 -3652
rect 321 -3800 331 -3640
rect 383 -3800 393 -3640
rect 430 -3652 476 -3640
rect 142 -4040 188 -4028
rect 225 -4040 235 -3880
rect 287 -4040 297 -3880
rect 334 -4028 340 -3800
rect 374 -4028 380 -3800
rect 430 -3880 436 -3652
rect 470 -3880 476 -3652
rect 513 -3800 523 -3640
rect 575 -3800 585 -3640
rect 622 -3652 668 -3640
rect 334 -4040 380 -4028
rect 417 -4040 427 -3880
rect 479 -4040 489 -3880
rect 526 -4028 532 -3800
rect 566 -4028 572 -3800
rect 622 -3880 628 -3652
rect 662 -3880 668 -3652
rect 705 -3800 715 -3640
rect 767 -3800 777 -3640
rect 814 -3652 860 -3640
rect 526 -4040 572 -4028
rect 609 -4040 619 -3880
rect 671 -4040 681 -3880
rect 718 -4028 724 -3800
rect 758 -4028 764 -3800
rect 814 -3880 820 -3652
rect 854 -3880 860 -3652
rect 897 -3800 907 -3640
rect 959 -3800 969 -3640
rect 1006 -3652 1052 -3640
rect 718 -4040 764 -4028
rect 801 -4040 811 -3880
rect 863 -4040 873 -3880
rect 910 -4028 916 -3800
rect 950 -4028 956 -3800
rect 1006 -3880 1012 -3652
rect 1046 -3880 1052 -3652
rect 1089 -3800 1099 -3640
rect 1151 -3800 1161 -3640
rect 1198 -3652 1244 -3640
rect 910 -4040 956 -4028
rect 993 -4040 1003 -3880
rect 1055 -4040 1065 -3880
rect 1102 -4028 1108 -3800
rect 1142 -4028 1148 -3800
rect 1198 -3880 1204 -3652
rect 1238 -3880 1244 -3652
rect 1102 -4040 1148 -4028
rect 1185 -4040 1195 -3880
rect 1247 -4040 1257 -3880
rect -1160 -4077 -1102 -4072
rect -968 -4077 -910 -4072
rect -776 -4077 -718 -4072
rect -584 -4077 -526 -4072
rect -392 -4077 -334 -4072
rect -200 -4077 -142 -4072
rect -8 -4077 50 -4072
rect 184 -4077 242 -4072
rect 376 -4077 434 -4072
rect 568 -4077 626 -4072
rect 760 -4077 818 -4072
rect 952 -4077 1010 -4072
rect 1144 -4077 1202 -4072
rect -1203 -4078 1247 -4077
rect -1203 -4080 -1148 -4078
rect -1270 -4112 -1148 -4080
rect -1114 -4112 -956 -4078
rect -922 -4112 -764 -4078
rect -730 -4112 -572 -4078
rect -538 -4112 -380 -4078
rect -346 -4112 -188 -4078
rect -154 -4112 4 -4078
rect 38 -4112 196 -4078
rect 230 -4112 388 -4078
rect 422 -4112 580 -4078
rect 614 -4112 772 -4078
rect 806 -4112 964 -4078
rect 998 -4112 1156 -4078
rect 1190 -4112 1247 -4078
rect -1270 -4120 1247 -4112
rect -1346 -4127 1247 -4120
rect -1346 -4130 -1196 -4127
rect -1386 -4428 -1136 -4420
rect 284 -4428 674 -4420
rect -1386 -4444 2093 -4428
rect -1386 -4478 -1127 -4444
rect -1093 -4478 -1029 -4444
rect -995 -4478 -931 -4444
rect -897 -4478 -833 -4444
rect -799 -4478 -735 -4444
rect -701 -4478 -637 -4444
rect -603 -4478 -539 -4444
rect -505 -4478 -441 -4444
rect -407 -4478 -343 -4444
rect -309 -4478 -245 -4444
rect -211 -4478 -147 -4444
rect -113 -4478 -49 -4444
rect -15 -4478 49 -4444
rect 83 -4478 147 -4444
rect 181 -4478 245 -4444
rect 279 -4478 671 -4444
rect 705 -4478 769 -4444
rect 803 -4478 867 -4444
rect 901 -4478 965 -4444
rect 999 -4478 1063 -4444
rect 1097 -4478 1161 -4444
rect 1195 -4478 1259 -4444
rect 1293 -4478 1357 -4444
rect 1391 -4478 1455 -4444
rect 1489 -4478 1553 -4444
rect 1587 -4478 1651 -4444
rect 1685 -4478 1749 -4444
rect 1783 -4478 1847 -4444
rect 1881 -4478 1945 -4444
rect 1979 -4478 2043 -4444
rect 2077 -4478 2093 -4444
rect -1386 -4490 2093 -4478
rect -1386 -4960 -1236 -4490
rect -1143 -4494 295 -4490
rect -1182 -4537 -1136 -4525
rect -1182 -4765 -1176 -4537
rect -1142 -4765 -1136 -4537
rect -1097 -4685 -1087 -4525
rect -1035 -4685 -1025 -4525
rect -986 -4537 -940 -4525
rect -1195 -4925 -1185 -4765
rect -1133 -4925 -1123 -4765
rect -1084 -4913 -1078 -4685
rect -1044 -4913 -1038 -4685
rect -986 -4765 -980 -4537
rect -946 -4765 -940 -4537
rect -901 -4685 -891 -4525
rect -839 -4685 -829 -4525
rect -790 -4537 -744 -4525
rect -1084 -4925 -1038 -4913
rect -999 -4925 -989 -4765
rect -937 -4925 -927 -4765
rect -888 -4913 -882 -4685
rect -848 -4913 -842 -4685
rect -790 -4765 -784 -4537
rect -750 -4765 -744 -4537
rect -705 -4685 -695 -4525
rect -643 -4685 -633 -4525
rect -594 -4537 -548 -4525
rect -888 -4925 -842 -4913
rect -803 -4925 -793 -4765
rect -741 -4925 -731 -4765
rect -692 -4913 -686 -4685
rect -652 -4913 -646 -4685
rect -594 -4765 -588 -4537
rect -554 -4765 -548 -4537
rect -509 -4685 -499 -4525
rect -447 -4685 -437 -4525
rect -398 -4537 -352 -4525
rect -692 -4925 -646 -4913
rect -607 -4925 -597 -4765
rect -545 -4925 -535 -4765
rect -496 -4913 -490 -4685
rect -456 -4913 -450 -4685
rect -398 -4765 -392 -4537
rect -358 -4765 -352 -4537
rect -313 -4685 -303 -4525
rect -251 -4685 -241 -4525
rect -202 -4537 -156 -4525
rect -496 -4925 -450 -4913
rect -411 -4925 -401 -4765
rect -349 -4925 -339 -4765
rect -300 -4913 -294 -4685
rect -260 -4913 -254 -4685
rect -202 -4765 -196 -4537
rect -162 -4765 -156 -4537
rect -117 -4685 -107 -4525
rect -55 -4685 -45 -4525
rect -6 -4537 40 -4525
rect -300 -4925 -254 -4913
rect -215 -4925 -205 -4765
rect -153 -4925 -143 -4765
rect -104 -4913 -98 -4685
rect -64 -4913 -58 -4685
rect -6 -4765 0 -4537
rect 34 -4765 40 -4537
rect 79 -4685 89 -4525
rect 141 -4685 151 -4525
rect 190 -4537 236 -4525
rect -104 -4925 -58 -4913
rect -19 -4925 -9 -4765
rect 43 -4925 53 -4765
rect 92 -4913 98 -4685
rect 132 -4913 138 -4685
rect 190 -4765 196 -4537
rect 230 -4765 236 -4537
rect 275 -4685 285 -4525
rect 337 -4685 347 -4525
rect 92 -4925 138 -4913
rect 177 -4925 187 -4765
rect 239 -4925 249 -4765
rect 288 -4913 294 -4685
rect 328 -4913 334 -4685
rect 288 -4925 334 -4913
rect -1143 -4960 295 -4956
rect 434 -4960 514 -4490
rect 655 -4494 2093 -4490
rect 616 -4537 662 -4525
rect 616 -4765 622 -4537
rect 656 -4765 662 -4537
rect 701 -4685 711 -4525
rect 763 -4685 773 -4525
rect 812 -4537 858 -4525
rect 603 -4925 613 -4765
rect 665 -4925 675 -4765
rect 714 -4913 720 -4685
rect 754 -4913 760 -4685
rect 812 -4765 818 -4537
rect 852 -4765 858 -4537
rect 897 -4685 907 -4525
rect 959 -4685 969 -4525
rect 1008 -4537 1054 -4525
rect 714 -4925 760 -4913
rect 799 -4925 809 -4765
rect 861 -4925 871 -4765
rect 910 -4913 916 -4685
rect 950 -4913 956 -4685
rect 1008 -4765 1014 -4537
rect 1048 -4765 1054 -4537
rect 1093 -4685 1103 -4525
rect 1155 -4685 1165 -4525
rect 1204 -4537 1250 -4525
rect 910 -4925 956 -4913
rect 995 -4925 1005 -4765
rect 1057 -4925 1067 -4765
rect 1106 -4913 1112 -4685
rect 1146 -4913 1152 -4685
rect 1204 -4765 1210 -4537
rect 1244 -4765 1250 -4537
rect 1289 -4685 1299 -4525
rect 1351 -4685 1361 -4525
rect 1400 -4537 1446 -4525
rect 1106 -4925 1152 -4913
rect 1191 -4925 1201 -4765
rect 1253 -4925 1263 -4765
rect 1302 -4913 1308 -4685
rect 1342 -4913 1348 -4685
rect 1400 -4765 1406 -4537
rect 1440 -4765 1446 -4537
rect 1485 -4685 1495 -4525
rect 1547 -4685 1557 -4525
rect 1596 -4537 1642 -4525
rect 1302 -4925 1348 -4913
rect 1387 -4925 1397 -4765
rect 1449 -4925 1459 -4765
rect 1498 -4913 1504 -4685
rect 1538 -4913 1544 -4685
rect 1596 -4765 1602 -4537
rect 1636 -4765 1642 -4537
rect 1681 -4685 1691 -4525
rect 1743 -4685 1753 -4525
rect 1792 -4537 1838 -4525
rect 1498 -4925 1544 -4913
rect 1583 -4925 1593 -4765
rect 1645 -4925 1655 -4765
rect 1694 -4913 1700 -4685
rect 1734 -4913 1740 -4685
rect 1792 -4765 1798 -4537
rect 1832 -4765 1838 -4537
rect 1877 -4685 1887 -4525
rect 1939 -4685 1949 -4525
rect 1988 -4537 2034 -4525
rect 1694 -4925 1740 -4913
rect 1779 -4925 1789 -4765
rect 1841 -4925 1851 -4765
rect 1890 -4913 1896 -4685
rect 1930 -4913 1936 -4685
rect 1988 -4765 1994 -4537
rect 2028 -4765 2034 -4537
rect 2073 -4685 2083 -4525
rect 2135 -4685 2145 -4525
rect 1890 -4925 1936 -4913
rect 1975 -4925 1985 -4765
rect 2037 -4925 2047 -4765
rect 2086 -4913 2092 -4685
rect 2126 -4913 2132 -4685
rect 2086 -4925 2132 -4913
rect 655 -4960 2093 -4956
rect -1386 -4972 2104 -4960
rect -1386 -5006 -1127 -4972
rect -1093 -5006 -1029 -4972
rect -995 -5006 -931 -4972
rect -897 -5006 -833 -4972
rect -799 -5006 -735 -4972
rect -701 -5006 -637 -4972
rect -603 -5006 -539 -4972
rect -505 -5006 -441 -4972
rect -407 -5006 -343 -4972
rect -309 -5006 -245 -4972
rect -211 -5006 -147 -4972
rect -113 -5006 -49 -4972
rect -15 -5006 49 -4972
rect 83 -5006 147 -4972
rect 181 -5006 245 -4972
rect 279 -5006 671 -4972
rect 705 -5006 769 -4972
rect 803 -5006 867 -4972
rect 901 -5006 965 -4972
rect 999 -5006 1063 -4972
rect 1097 -5006 1161 -4972
rect 1195 -5006 1259 -4972
rect 1293 -5006 1357 -4972
rect 1391 -5006 1455 -4972
rect 1489 -5006 1553 -4972
rect 1587 -5006 1651 -4972
rect 1685 -5006 1749 -4972
rect 1783 -5006 1847 -4972
rect 1881 -5006 1945 -4972
rect 1979 -5006 2043 -4972
rect 2077 -5006 2104 -4972
rect 2208 -5000 2350 -4988
rect -1386 -5080 2104 -5006
rect -1386 -5114 -1127 -5080
rect -1093 -5114 -1029 -5080
rect -995 -5114 -931 -5080
rect -897 -5114 -833 -5080
rect -799 -5114 -735 -5080
rect -701 -5114 -637 -5080
rect -603 -5114 -539 -5080
rect -505 -5114 -441 -5080
rect -407 -5114 -343 -5080
rect -309 -5114 -245 -5080
rect -211 -5114 -147 -5080
rect -113 -5114 -49 -5080
rect -15 -5114 49 -5080
rect 83 -5114 147 -5080
rect 181 -5114 245 -5080
rect 279 -5114 671 -5080
rect 705 -5114 769 -5080
rect 803 -5114 867 -5080
rect 901 -5114 965 -5080
rect 999 -5114 1063 -5080
rect 1097 -5114 1161 -5080
rect 1195 -5114 1259 -5080
rect 1293 -5114 1357 -5080
rect 1391 -5114 1455 -5080
rect 1489 -5114 1553 -5080
rect 1587 -5114 1651 -5080
rect 1685 -5114 1749 -5080
rect 1783 -5114 1847 -5080
rect 1881 -5114 1945 -5080
rect 1979 -5114 2043 -5080
rect 2077 -5114 2104 -5080
rect -1386 -5130 2104 -5114
rect -1386 -5600 -1236 -5130
rect -1195 -5321 -1185 -5161
rect -1133 -5321 -1123 -5161
rect -1084 -5173 -1038 -5161
rect -1182 -5549 -1176 -5321
rect -1142 -5549 -1136 -5321
rect -1084 -5401 -1078 -5173
rect -1044 -5401 -1038 -5173
rect -999 -5321 -989 -5161
rect -937 -5321 -927 -5161
rect -888 -5173 -842 -5161
rect -1182 -5561 -1136 -5549
rect -1097 -5561 -1087 -5401
rect -1035 -5561 -1025 -5401
rect -986 -5549 -980 -5321
rect -946 -5549 -940 -5321
rect -888 -5401 -882 -5173
rect -848 -5401 -842 -5173
rect -803 -5321 -793 -5161
rect -741 -5321 -731 -5161
rect -692 -5173 -646 -5161
rect -986 -5561 -940 -5549
rect -901 -5561 -891 -5401
rect -839 -5561 -829 -5401
rect -790 -5549 -784 -5321
rect -750 -5549 -744 -5321
rect -692 -5401 -686 -5173
rect -652 -5401 -646 -5173
rect -607 -5321 -597 -5161
rect -545 -5321 -535 -5161
rect -496 -5173 -450 -5161
rect -790 -5561 -744 -5549
rect -705 -5561 -695 -5401
rect -643 -5561 -633 -5401
rect -594 -5549 -588 -5321
rect -554 -5549 -548 -5321
rect -496 -5401 -490 -5173
rect -456 -5401 -450 -5173
rect -411 -5321 -401 -5161
rect -349 -5321 -339 -5161
rect -300 -5173 -254 -5161
rect -594 -5561 -548 -5549
rect -509 -5561 -499 -5401
rect -447 -5561 -437 -5401
rect -398 -5549 -392 -5321
rect -358 -5549 -352 -5321
rect -300 -5401 -294 -5173
rect -260 -5401 -254 -5173
rect -215 -5321 -205 -5161
rect -153 -5321 -143 -5161
rect -104 -5173 -58 -5161
rect -398 -5561 -352 -5549
rect -313 -5561 -303 -5401
rect -251 -5561 -241 -5401
rect -202 -5549 -196 -5321
rect -162 -5549 -156 -5321
rect -104 -5401 -98 -5173
rect -64 -5401 -58 -5173
rect -19 -5321 -9 -5161
rect 43 -5321 53 -5161
rect 92 -5173 138 -5161
rect -202 -5561 -156 -5549
rect -117 -5561 -107 -5401
rect -55 -5561 -45 -5401
rect -6 -5549 0 -5321
rect 34 -5549 40 -5321
rect 92 -5401 98 -5173
rect 132 -5401 138 -5173
rect 177 -5321 187 -5161
rect 239 -5321 249 -5161
rect 288 -5173 334 -5161
rect -6 -5561 40 -5549
rect 79 -5561 89 -5401
rect 141 -5561 151 -5401
rect 190 -5549 196 -5321
rect 230 -5549 236 -5321
rect 288 -5401 294 -5173
rect 328 -5401 334 -5173
rect 190 -5561 236 -5549
rect 275 -5561 285 -5401
rect 337 -5561 347 -5401
rect 434 -5590 514 -5130
rect 603 -5321 613 -5161
rect 665 -5321 675 -5161
rect 714 -5173 760 -5161
rect 616 -5549 622 -5321
rect 656 -5549 662 -5321
rect 714 -5401 720 -5173
rect 754 -5401 760 -5173
rect 799 -5321 809 -5161
rect 861 -5321 871 -5161
rect 910 -5173 956 -5161
rect 616 -5561 662 -5549
rect 701 -5561 711 -5401
rect 763 -5561 773 -5401
rect 812 -5549 818 -5321
rect 852 -5549 858 -5321
rect 910 -5401 916 -5173
rect 950 -5401 956 -5173
rect 995 -5321 1005 -5161
rect 1057 -5321 1067 -5161
rect 1106 -5173 1152 -5161
rect 812 -5561 858 -5549
rect 897 -5561 907 -5401
rect 959 -5561 969 -5401
rect 1008 -5549 1014 -5321
rect 1048 -5549 1054 -5321
rect 1106 -5401 1112 -5173
rect 1146 -5401 1152 -5173
rect 1191 -5321 1201 -5161
rect 1253 -5321 1263 -5161
rect 1302 -5173 1348 -5161
rect 1008 -5561 1054 -5549
rect 1093 -5561 1103 -5401
rect 1155 -5561 1165 -5401
rect 1204 -5549 1210 -5321
rect 1244 -5549 1250 -5321
rect 1302 -5401 1308 -5173
rect 1342 -5401 1348 -5173
rect 1387 -5321 1397 -5161
rect 1449 -5321 1459 -5161
rect 1498 -5173 1544 -5161
rect 1204 -5561 1250 -5549
rect 1289 -5561 1299 -5401
rect 1351 -5561 1361 -5401
rect 1400 -5549 1406 -5321
rect 1440 -5549 1446 -5321
rect 1498 -5401 1504 -5173
rect 1538 -5401 1544 -5173
rect 1583 -5321 1593 -5161
rect 1645 -5321 1655 -5161
rect 1694 -5173 1740 -5161
rect 1400 -5561 1446 -5549
rect 1485 -5561 1495 -5401
rect 1547 -5561 1557 -5401
rect 1596 -5549 1602 -5321
rect 1636 -5549 1642 -5321
rect 1694 -5401 1700 -5173
rect 1734 -5401 1740 -5173
rect 1779 -5321 1789 -5161
rect 1841 -5321 1851 -5161
rect 1890 -5173 1936 -5161
rect 1596 -5561 1642 -5549
rect 1681 -5561 1691 -5401
rect 1743 -5561 1753 -5401
rect 1792 -5549 1798 -5321
rect 1832 -5549 1838 -5321
rect 1890 -5401 1896 -5173
rect 1930 -5401 1936 -5173
rect 1975 -5321 1985 -5161
rect 2037 -5321 2047 -5161
rect 2086 -5173 2132 -5161
rect 1792 -5561 1838 -5549
rect 1877 -5561 1887 -5401
rect 1939 -5561 1949 -5401
rect 1988 -5549 1994 -5321
rect 2028 -5549 2034 -5321
rect 2086 -5401 2092 -5173
rect 2126 -5401 2132 -5173
rect 1988 -5561 2034 -5549
rect 2073 -5561 2083 -5401
rect 2135 -5561 2145 -5401
rect 2204 -5560 2214 -5000
rect 2344 -5560 2354 -5000
rect 4180 -5090 4190 -5080
rect 2474 -5096 4190 -5090
rect 2474 -5130 2486 -5096
rect 2554 -5130 2644 -5096
rect 2712 -5130 2802 -5096
rect 2870 -5130 2960 -5096
rect 3028 -5130 3118 -5096
rect 3186 -5130 3276 -5096
rect 3344 -5130 3434 -5096
rect 3502 -5130 3592 -5096
rect 3660 -5130 3750 -5096
rect 3818 -5130 3908 -5096
rect 3976 -5130 4190 -5096
rect 2474 -5136 2566 -5130
rect 2632 -5136 2724 -5130
rect 2790 -5136 2882 -5130
rect 2948 -5136 3040 -5130
rect 3106 -5136 3198 -5130
rect 3264 -5136 3356 -5130
rect 3422 -5136 3514 -5130
rect 3580 -5136 3672 -5130
rect 3738 -5136 3830 -5130
rect 3896 -5136 3988 -5130
rect 2418 -5189 2464 -5177
rect 2418 -5417 2424 -5189
rect 2458 -5417 2464 -5189
rect 2563 -5337 2573 -5177
rect 2625 -5337 2635 -5177
rect 2734 -5189 2780 -5177
rect 2208 -5572 2350 -5560
rect 2405 -5577 2415 -5417
rect 2467 -5577 2477 -5417
rect 2576 -5565 2582 -5337
rect 2616 -5565 2622 -5337
rect 2734 -5417 2740 -5189
rect 2774 -5417 2780 -5189
rect 2879 -5337 2889 -5177
rect 2941 -5337 2951 -5177
rect 3050 -5189 3096 -5177
rect 2576 -5577 2622 -5565
rect 2721 -5577 2731 -5417
rect 2783 -5577 2793 -5417
rect 2892 -5565 2898 -5337
rect 2932 -5565 2938 -5337
rect 3050 -5417 3056 -5189
rect 3090 -5417 3096 -5189
rect 3195 -5337 3205 -5177
rect 3257 -5337 3267 -5177
rect 3366 -5189 3412 -5177
rect 2892 -5577 2938 -5565
rect 3037 -5577 3047 -5417
rect 3099 -5577 3109 -5417
rect 3208 -5565 3214 -5337
rect 3248 -5565 3254 -5337
rect 3366 -5417 3372 -5189
rect 3406 -5417 3412 -5189
rect 3511 -5337 3521 -5177
rect 3573 -5337 3583 -5177
rect 3682 -5189 3728 -5177
rect 3208 -5577 3254 -5565
rect 3353 -5577 3363 -5417
rect 3415 -5577 3425 -5417
rect 3524 -5565 3530 -5337
rect 3564 -5565 3570 -5337
rect 3682 -5417 3688 -5189
rect 3722 -5417 3728 -5189
rect 3827 -5337 3837 -5177
rect 3889 -5337 3899 -5177
rect 3998 -5189 4044 -5177
rect 3524 -5577 3570 -5565
rect 3669 -5577 3679 -5417
rect 3731 -5577 3741 -5417
rect 3840 -5565 3846 -5337
rect 3880 -5565 3886 -5337
rect 3998 -5417 4004 -5189
rect 4038 -5417 4044 -5189
rect 4090 -5190 4190 -5130
rect 3840 -5577 3886 -5565
rect 3985 -5577 3995 -5417
rect 4047 -5577 4057 -5417
rect 284 -5592 674 -5590
rect -1143 -5600 2093 -5592
rect -1386 -5608 2093 -5600
rect -1386 -5642 -1127 -5608
rect -1093 -5642 -1029 -5608
rect -995 -5642 -931 -5608
rect -897 -5642 -833 -5608
rect -799 -5642 -735 -5608
rect -701 -5642 -637 -5608
rect -603 -5642 -539 -5608
rect -505 -5642 -441 -5608
rect -407 -5642 -343 -5608
rect -309 -5642 -245 -5608
rect -211 -5642 -147 -5608
rect -113 -5642 -49 -5608
rect -15 -5642 49 -5608
rect 83 -5642 147 -5608
rect 181 -5642 245 -5608
rect 279 -5642 671 -5608
rect 705 -5642 769 -5608
rect 803 -5642 867 -5608
rect 901 -5642 965 -5608
rect 999 -5642 1063 -5608
rect 1097 -5642 1161 -5608
rect 1195 -5642 1259 -5608
rect 1293 -5642 1357 -5608
rect 1391 -5642 1455 -5608
rect 1489 -5642 1553 -5608
rect 1587 -5642 1651 -5608
rect 1685 -5642 1749 -5608
rect 1783 -5642 1847 -5608
rect 1881 -5642 1945 -5608
rect 1979 -5642 2043 -5608
rect 2077 -5642 2093 -5608
rect 2474 -5624 2566 -5618
rect 2474 -5630 2486 -5624
rect -1386 -5658 2093 -5642
rect 2464 -5658 2486 -5630
rect 2554 -5630 2566 -5624
rect 2632 -5624 2724 -5618
rect 2632 -5630 2644 -5624
rect 2554 -5658 2644 -5630
rect 2712 -5630 2724 -5624
rect 2790 -5624 2882 -5618
rect 2790 -5630 2802 -5624
rect 2712 -5658 2802 -5630
rect 2870 -5630 2882 -5624
rect 2948 -5624 3040 -5618
rect 2948 -5630 2960 -5624
rect 2870 -5658 2960 -5630
rect 3028 -5630 3040 -5624
rect 3106 -5624 3198 -5618
rect 3106 -5630 3118 -5624
rect 3028 -5658 3118 -5630
rect 3186 -5630 3198 -5624
rect 3264 -5624 3356 -5618
rect 3264 -5630 3276 -5624
rect 3186 -5658 3276 -5630
rect 3344 -5630 3356 -5624
rect 3422 -5624 3514 -5618
rect 3422 -5630 3434 -5624
rect 3344 -5658 3434 -5630
rect 3502 -5630 3514 -5624
rect 3580 -5624 3672 -5618
rect 3580 -5630 3592 -5624
rect 3502 -5658 3592 -5630
rect 3660 -5630 3672 -5624
rect 3738 -5624 3830 -5618
rect 3738 -5630 3750 -5624
rect 3660 -5658 3750 -5630
rect 3818 -5630 3830 -5624
rect 3896 -5624 3988 -5618
rect 3896 -5630 3908 -5624
rect 3818 -5658 3908 -5630
rect 3976 -5630 3988 -5624
rect 4094 -5630 4134 -5190
rect 4180 -5200 4190 -5190
rect 4290 -5200 4300 -5080
rect 3976 -5658 4134 -5630
rect -1386 -5670 -1136 -5658
rect 284 -5660 674 -5658
rect -1386 -5890 -1236 -5670
rect 434 -5850 514 -5660
rect 2464 -5670 4134 -5658
rect -1386 -5904 -1136 -5890
rect 434 -5904 1544 -5850
rect -1386 -5920 1544 -5904
rect -1386 -5954 -1127 -5920
rect -1093 -5954 -1030 -5920
rect -996 -5954 -931 -5920
rect -897 -5954 -834 -5920
rect -800 -5954 -735 -5920
rect -701 -5954 -638 -5920
rect -604 -5954 -539 -5920
rect -505 -5954 -442 -5920
rect -408 -5954 -343 -5920
rect -309 -5954 -246 -5920
rect -212 -5954 -147 -5920
rect -113 -5954 -50 -5920
rect -16 -5954 49 -5920
rect 83 -5954 146 -5920
rect 180 -5954 245 -5920
rect 279 -5954 342 -5920
rect 376 -5954 441 -5920
rect 475 -5954 538 -5920
rect 572 -5954 637 -5920
rect 671 -5954 734 -5920
rect 768 -5954 833 -5920
rect 867 -5954 930 -5920
rect 964 -5954 1029 -5920
rect 1063 -5954 1126 -5920
rect 1160 -5954 1225 -5920
rect 1259 -5954 1544 -5920
rect -1386 -5960 1544 -5954
rect -1386 -6430 -1236 -5960
rect -1144 -5964 1274 -5960
rect -1182 -6004 -1136 -5992
rect -1182 -6232 -1176 -6004
rect -1142 -6232 -1136 -6004
rect -1097 -6152 -1087 -5992
rect -1035 -6152 -1025 -5992
rect -986 -6004 -940 -5992
rect -1195 -6392 -1185 -6232
rect -1133 -6392 -1123 -6232
rect -1084 -6380 -1078 -6152
rect -1044 -6380 -1038 -6152
rect -986 -6232 -980 -6004
rect -946 -6232 -940 -6004
rect -901 -6152 -891 -5992
rect -839 -6152 -829 -5992
rect -790 -6004 -744 -5992
rect -1084 -6392 -1038 -6380
rect -999 -6392 -989 -6232
rect -937 -6392 -927 -6232
rect -888 -6380 -882 -6152
rect -848 -6380 -842 -6152
rect -790 -6232 -784 -6004
rect -750 -6232 -744 -6004
rect -705 -6152 -695 -5992
rect -643 -6152 -633 -5992
rect -594 -6004 -548 -5992
rect -888 -6392 -842 -6380
rect -803 -6392 -793 -6232
rect -741 -6392 -731 -6232
rect -692 -6380 -686 -6152
rect -652 -6380 -646 -6152
rect -594 -6232 -588 -6004
rect -554 -6232 -548 -6004
rect -509 -6152 -499 -5992
rect -447 -6152 -437 -5992
rect -398 -6004 -352 -5992
rect -692 -6392 -646 -6380
rect -607 -6392 -597 -6232
rect -545 -6392 -535 -6232
rect -496 -6380 -490 -6152
rect -456 -6380 -450 -6152
rect -398 -6232 -392 -6004
rect -358 -6232 -352 -6004
rect -313 -6152 -303 -5992
rect -251 -6152 -241 -5992
rect -202 -6004 -156 -5992
rect -496 -6392 -450 -6380
rect -411 -6392 -401 -6232
rect -349 -6392 -339 -6232
rect -300 -6380 -294 -6152
rect -260 -6380 -254 -6152
rect -202 -6232 -196 -6004
rect -162 -6232 -156 -6004
rect -117 -6152 -107 -5992
rect -55 -6152 -45 -5992
rect -6 -6004 40 -5992
rect -300 -6392 -254 -6380
rect -215 -6392 -205 -6232
rect -153 -6392 -143 -6232
rect -104 -6380 -98 -6152
rect -64 -6380 -58 -6152
rect -6 -6232 0 -6004
rect 34 -6232 40 -6004
rect 79 -6152 89 -5992
rect 141 -6152 151 -5992
rect 190 -6004 236 -5992
rect -104 -6392 -58 -6380
rect -19 -6392 -9 -6232
rect 43 -6392 53 -6232
rect 92 -6380 98 -6152
rect 132 -6380 138 -6152
rect 190 -6232 196 -6004
rect 230 -6232 236 -6004
rect 275 -6152 285 -5992
rect 337 -6152 347 -5992
rect 386 -6004 432 -5992
rect 92 -6392 138 -6380
rect 177 -6392 187 -6232
rect 239 -6392 249 -6232
rect 288 -6380 294 -6152
rect 328 -6380 334 -6152
rect 386 -6232 392 -6004
rect 426 -6232 432 -6004
rect 471 -6152 481 -5992
rect 533 -6152 543 -5992
rect 582 -6004 628 -5992
rect 288 -6392 334 -6380
rect 373 -6392 383 -6232
rect 435 -6392 445 -6232
rect 484 -6380 490 -6152
rect 524 -6380 530 -6152
rect 582 -6232 588 -6004
rect 622 -6232 628 -6004
rect 667 -6152 677 -5992
rect 729 -6152 739 -5992
rect 778 -6004 824 -5992
rect 484 -6392 530 -6380
rect 569 -6392 579 -6232
rect 631 -6392 641 -6232
rect 680 -6380 686 -6152
rect 720 -6380 726 -6152
rect 778 -6232 784 -6004
rect 818 -6232 824 -6004
rect 863 -6152 873 -5992
rect 925 -6152 935 -5992
rect 974 -6004 1020 -5992
rect 680 -6392 726 -6380
rect 765 -6392 775 -6232
rect 827 -6392 837 -6232
rect 876 -6380 882 -6152
rect 916 -6380 922 -6152
rect 974 -6232 980 -6004
rect 1014 -6232 1020 -6004
rect 1059 -6152 1069 -5992
rect 1121 -6152 1131 -5992
rect 1170 -6004 1216 -5992
rect 876 -6392 922 -6380
rect 961 -6392 971 -6232
rect 1023 -6392 1033 -6232
rect 1072 -6380 1078 -6152
rect 1112 -6380 1118 -6152
rect 1170 -6232 1176 -6004
rect 1210 -6232 1216 -6004
rect 1255 -6152 1265 -5992
rect 1317 -6152 1327 -5992
rect 1072 -6392 1118 -6380
rect 1157 -6392 1167 -6232
rect 1219 -6392 1229 -6232
rect 1268 -6380 1274 -6152
rect 1308 -6380 1314 -6152
rect 1268 -6392 1314 -6380
rect -1144 -6430 1274 -6420
rect 1404 -6430 1544 -5960
rect 2154 -6410 2164 -6220
rect 2414 -6224 3954 -6220
rect 2414 -6240 3955 -6224
rect 2414 -6274 2533 -6240
rect 2567 -6274 2631 -6240
rect 2665 -6274 2729 -6240
rect 2763 -6274 2827 -6240
rect 2861 -6274 2925 -6240
rect 2959 -6274 3023 -6240
rect 3057 -6274 3121 -6240
rect 3155 -6274 3219 -6240
rect 3253 -6274 3317 -6240
rect 3351 -6274 3415 -6240
rect 3449 -6274 3513 -6240
rect 3547 -6274 3611 -6240
rect 3645 -6274 3709 -6240
rect 3743 -6274 3807 -6240
rect 3841 -6274 3905 -6240
rect 3939 -6274 3955 -6240
rect 2414 -6280 3955 -6274
rect 2414 -6410 2434 -6280
rect -1386 -6464 -1128 -6430
rect -1094 -6464 -1029 -6430
rect -995 -6464 -932 -6430
rect -898 -6464 -833 -6430
rect -799 -6464 -736 -6430
rect -702 -6464 -637 -6430
rect -603 -6464 -540 -6430
rect -506 -6464 -441 -6430
rect -407 -6464 -344 -6430
rect -310 -6464 -245 -6430
rect -211 -6464 -148 -6430
rect -114 -6464 -49 -6430
rect -15 -6464 48 -6430
rect 82 -6464 147 -6430
rect 181 -6464 244 -6430
rect 278 -6464 343 -6430
rect 377 -6464 440 -6430
rect 474 -6464 539 -6430
rect 573 -6464 636 -6430
rect 670 -6464 735 -6430
rect 769 -6464 832 -6430
rect 866 -6464 931 -6430
rect 965 -6464 1028 -6430
rect 1062 -6464 1127 -6430
rect 1161 -6464 1224 -6430
rect 1258 -6464 1544 -6430
rect -1386 -6538 1544 -6464
rect -1386 -6572 -1127 -6538
rect -1093 -6572 -1029 -6538
rect -995 -6572 -931 -6538
rect -897 -6572 -833 -6538
rect -799 -6572 -735 -6538
rect -701 -6572 -637 -6538
rect -603 -6572 -539 -6538
rect -505 -6572 -441 -6538
rect -407 -6572 -343 -6538
rect -309 -6572 -245 -6538
rect -211 -6572 -147 -6538
rect -113 -6572 -49 -6538
rect -15 -6572 49 -6538
rect 83 -6572 147 -6538
rect 181 -6572 245 -6538
rect 279 -6572 343 -6538
rect 377 -6572 441 -6538
rect 475 -6572 539 -6538
rect 573 -6572 637 -6538
rect 671 -6572 735 -6538
rect 769 -6572 833 -6538
rect 867 -6572 931 -6538
rect 965 -6572 1029 -6538
rect 1063 -6572 1127 -6538
rect 1161 -6572 1225 -6538
rect 1259 -6572 1544 -6538
rect -1386 -6580 1544 -6572
rect -1386 -7040 -1236 -6580
rect -1143 -6582 1275 -6580
rect -1195 -6770 -1185 -6610
rect -1133 -6770 -1123 -6610
rect -1084 -6622 -1038 -6610
rect -1182 -6998 -1176 -6770
rect -1142 -6998 -1136 -6770
rect -1084 -6850 -1078 -6622
rect -1044 -6850 -1038 -6622
rect -999 -6770 -989 -6610
rect -937 -6770 -927 -6610
rect -888 -6622 -842 -6610
rect -1182 -7010 -1136 -6998
rect -1097 -7010 -1087 -6850
rect -1035 -7010 -1025 -6850
rect -986 -6998 -980 -6770
rect -946 -6998 -940 -6770
rect -888 -6850 -882 -6622
rect -848 -6850 -842 -6622
rect -803 -6770 -793 -6610
rect -741 -6770 -731 -6610
rect -692 -6622 -646 -6610
rect -986 -7010 -940 -6998
rect -901 -7010 -891 -6850
rect -839 -7010 -829 -6850
rect -790 -6998 -784 -6770
rect -750 -6998 -744 -6770
rect -692 -6850 -686 -6622
rect -652 -6850 -646 -6622
rect -607 -6770 -597 -6610
rect -545 -6770 -535 -6610
rect -496 -6622 -450 -6610
rect -790 -7010 -744 -6998
rect -705 -7010 -695 -6850
rect -643 -7010 -633 -6850
rect -594 -6998 -588 -6770
rect -554 -6998 -548 -6770
rect -496 -6850 -490 -6622
rect -456 -6850 -450 -6622
rect -411 -6770 -401 -6610
rect -349 -6770 -339 -6610
rect -300 -6622 -254 -6610
rect -594 -7010 -548 -6998
rect -509 -7010 -499 -6850
rect -447 -7010 -437 -6850
rect -398 -6998 -392 -6770
rect -358 -6998 -352 -6770
rect -300 -6850 -294 -6622
rect -260 -6850 -254 -6622
rect -215 -6770 -205 -6610
rect -153 -6770 -143 -6610
rect -104 -6622 -58 -6610
rect -398 -7010 -352 -6998
rect -313 -7010 -303 -6850
rect -251 -7010 -241 -6850
rect -202 -6998 -196 -6770
rect -162 -6998 -156 -6770
rect -104 -6850 -98 -6622
rect -64 -6850 -58 -6622
rect -19 -6770 -9 -6610
rect 43 -6770 53 -6610
rect 92 -6622 138 -6610
rect -202 -7010 -156 -6998
rect -117 -7010 -107 -6850
rect -55 -7010 -45 -6850
rect -6 -6998 0 -6770
rect 34 -6998 40 -6770
rect 92 -6850 98 -6622
rect 132 -6850 138 -6622
rect 177 -6770 187 -6610
rect 239 -6770 249 -6610
rect 288 -6622 334 -6610
rect -6 -7010 40 -6998
rect 79 -7010 89 -6850
rect 141 -7010 151 -6850
rect 190 -6998 196 -6770
rect 230 -6998 236 -6770
rect 288 -6850 294 -6622
rect 328 -6850 334 -6622
rect 373 -6770 383 -6610
rect 435 -6770 445 -6610
rect 484 -6622 530 -6610
rect 190 -7010 236 -6998
rect 275 -7010 285 -6850
rect 337 -7010 347 -6850
rect 386 -6998 392 -6770
rect 426 -6998 432 -6770
rect 484 -6850 490 -6622
rect 524 -6850 530 -6622
rect 569 -6770 579 -6610
rect 631 -6770 641 -6610
rect 680 -6622 726 -6610
rect 386 -7010 432 -6998
rect 471 -7010 481 -6850
rect 533 -7010 543 -6850
rect 582 -6998 588 -6770
rect 622 -6998 628 -6770
rect 680 -6850 686 -6622
rect 720 -6850 726 -6622
rect 765 -6770 775 -6610
rect 827 -6770 837 -6610
rect 876 -6622 922 -6610
rect 582 -7010 628 -6998
rect 667 -7010 677 -6850
rect 729 -7010 739 -6850
rect 778 -6998 784 -6770
rect 818 -6998 824 -6770
rect 876 -6850 882 -6622
rect 916 -6850 922 -6622
rect 961 -6770 971 -6610
rect 1023 -6770 1033 -6610
rect 1072 -6622 1118 -6610
rect 778 -7010 824 -6998
rect 863 -7010 873 -6850
rect 925 -7010 935 -6850
rect 974 -6998 980 -6770
rect 1014 -6998 1020 -6770
rect 1072 -6850 1078 -6622
rect 1112 -6850 1118 -6622
rect 1157 -6770 1167 -6610
rect 1219 -6770 1229 -6610
rect 1268 -6622 1314 -6610
rect 974 -7010 1020 -6998
rect 1059 -7010 1069 -6850
rect 1121 -7010 1131 -6850
rect 1170 -6998 1176 -6770
rect 1210 -6998 1216 -6770
rect 1268 -6850 1274 -6622
rect 1308 -6850 1314 -6622
rect 1404 -6750 1544 -6580
rect 2198 -6750 2290 -6738
rect 2344 -6750 2434 -6410
rect 2465 -6472 2475 -6312
rect 2527 -6472 2537 -6312
rect 2576 -6324 2622 -6312
rect 2478 -6700 2484 -6472
rect 2518 -6700 2524 -6472
rect 2576 -6552 2582 -6324
rect 2616 -6552 2622 -6324
rect 2661 -6472 2671 -6312
rect 2723 -6472 2733 -6312
rect 2772 -6324 2818 -6312
rect 2478 -6712 2524 -6700
rect 2563 -6712 2573 -6552
rect 2625 -6712 2635 -6552
rect 2674 -6700 2680 -6472
rect 2714 -6700 2720 -6472
rect 2772 -6552 2778 -6324
rect 2812 -6552 2818 -6324
rect 2857 -6472 2867 -6312
rect 2919 -6472 2929 -6312
rect 2968 -6324 3014 -6312
rect 2674 -6712 2720 -6700
rect 2759 -6712 2769 -6552
rect 2821 -6712 2831 -6552
rect 2870 -6700 2876 -6472
rect 2910 -6700 2916 -6472
rect 2968 -6552 2974 -6324
rect 3008 -6552 3014 -6324
rect 3053 -6472 3063 -6312
rect 3115 -6472 3125 -6312
rect 3164 -6324 3210 -6312
rect 2870 -6712 2916 -6700
rect 2955 -6712 2965 -6552
rect 3017 -6712 3027 -6552
rect 3066 -6700 3072 -6472
rect 3106 -6700 3112 -6472
rect 3164 -6552 3170 -6324
rect 3204 -6552 3210 -6324
rect 3249 -6472 3259 -6312
rect 3311 -6472 3321 -6312
rect 3360 -6324 3406 -6312
rect 3066 -6712 3112 -6700
rect 3151 -6712 3161 -6552
rect 3213 -6712 3223 -6552
rect 3262 -6700 3268 -6472
rect 3302 -6700 3308 -6472
rect 3360 -6552 3366 -6324
rect 3400 -6552 3406 -6324
rect 3445 -6472 3455 -6312
rect 3507 -6472 3517 -6312
rect 3556 -6324 3602 -6312
rect 3262 -6712 3308 -6700
rect 3347 -6712 3357 -6552
rect 3409 -6712 3419 -6552
rect 3458 -6700 3464 -6472
rect 3498 -6700 3504 -6472
rect 3556 -6552 3562 -6324
rect 3596 -6552 3602 -6324
rect 3641 -6472 3651 -6312
rect 3703 -6472 3713 -6312
rect 3752 -6324 3798 -6312
rect 3458 -6712 3504 -6700
rect 3543 -6712 3553 -6552
rect 3605 -6712 3615 -6552
rect 3654 -6700 3660 -6472
rect 3694 -6700 3700 -6472
rect 3752 -6552 3758 -6324
rect 3792 -6552 3798 -6324
rect 3837 -6472 3847 -6312
rect 3899 -6472 3909 -6312
rect 3948 -6324 3994 -6312
rect 3654 -6712 3700 -6700
rect 3739 -6712 3749 -6552
rect 3801 -6712 3811 -6552
rect 3850 -6700 3856 -6472
rect 3890 -6700 3896 -6472
rect 3948 -6552 3954 -6324
rect 3988 -6552 3994 -6324
rect 3850 -6712 3896 -6700
rect 3935 -6712 3945 -6552
rect 3997 -6712 4007 -6552
rect 4048 -6730 4180 -6718
rect 2517 -6750 3955 -6744
rect 1170 -7010 1216 -6998
rect 1255 -7010 1265 -6850
rect 1317 -7010 1327 -6850
rect 1404 -6910 1454 -6750
rect 1684 -6910 1694 -6750
rect 2194 -6910 2204 -6750
rect 2284 -6910 2294 -6750
rect 2344 -6784 2533 -6750
rect 2567 -6784 2631 -6750
rect 2665 -6784 2729 -6750
rect 2763 -6784 2827 -6750
rect 2861 -6784 2925 -6750
rect 2959 -6784 3023 -6750
rect 3057 -6784 3121 -6750
rect 3155 -6784 3219 -6750
rect 3253 -6784 3317 -6750
rect 3351 -6784 3415 -6750
rect 3449 -6784 3513 -6750
rect 3547 -6784 3611 -6750
rect 3645 -6784 3709 -6750
rect 3743 -6784 3807 -6750
rect 3841 -6784 3905 -6750
rect 3939 -6784 3955 -6750
rect 2344 -6800 3955 -6784
rect 2344 -6842 3954 -6800
rect 2344 -6858 3955 -6842
rect 2344 -6890 2533 -6858
rect -1143 -7040 1275 -7038
rect 1404 -7040 1544 -6910
rect 2198 -6922 2290 -6910
rect -1386 -7048 1544 -7040
rect -1386 -7082 -1127 -7048
rect -1093 -7082 -1029 -7048
rect -995 -7082 -931 -7048
rect -897 -7082 -833 -7048
rect -799 -7082 -735 -7048
rect -701 -7082 -637 -7048
rect -603 -7082 -539 -7048
rect -505 -7082 -441 -7048
rect -407 -7082 -343 -7048
rect -309 -7082 -245 -7048
rect -211 -7082 -147 -7048
rect -113 -7082 -49 -7048
rect -15 -7082 49 -7048
rect 83 -7082 147 -7048
rect 181 -7082 245 -7048
rect 279 -7082 343 -7048
rect 377 -7082 441 -7048
rect 475 -7082 539 -7048
rect 573 -7082 637 -7048
rect 671 -7082 735 -7048
rect 769 -7082 833 -7048
rect 867 -7082 931 -7048
rect 965 -7082 1029 -7048
rect 1063 -7082 1127 -7048
rect 1161 -7082 1225 -7048
rect 1259 -7082 1544 -7048
rect -1386 -7098 1544 -7082
rect -1386 -7100 -1136 -7098
rect 1274 -7100 1544 -7098
rect -1386 -7330 -1236 -7100
rect -1386 -7348 -1136 -7330
rect 1404 -7340 1544 -7100
rect 1274 -7348 1544 -7340
rect -1386 -7364 1544 -7348
rect -1386 -7398 -1127 -7364
rect -1093 -7398 -1030 -7364
rect -996 -7398 -931 -7364
rect -897 -7398 -834 -7364
rect -800 -7398 -735 -7364
rect -701 -7398 -638 -7364
rect -604 -7398 -539 -7364
rect -505 -7398 -442 -7364
rect -408 -7398 -343 -7364
rect -309 -7398 -246 -7364
rect -212 -7398 -147 -7364
rect -113 -7398 -50 -7364
rect -16 -7398 49 -7364
rect 83 -7398 146 -7364
rect 180 -7398 245 -7364
rect 279 -7398 342 -7364
rect 376 -7398 441 -7364
rect 475 -7398 538 -7364
rect 572 -7398 637 -7364
rect 671 -7398 734 -7364
rect 768 -7398 833 -7364
rect 867 -7398 930 -7364
rect 964 -7398 1029 -7364
rect 1063 -7398 1126 -7364
rect 1160 -7398 1225 -7364
rect 1259 -7398 1544 -7364
rect -1386 -7400 1544 -7398
rect -1386 -7870 -1236 -7400
rect -1144 -7408 1274 -7400
rect -1182 -7448 -1136 -7436
rect -1182 -7676 -1176 -7448
rect -1142 -7676 -1136 -7448
rect -1097 -7596 -1087 -7436
rect -1035 -7596 -1025 -7436
rect -986 -7448 -940 -7436
rect -1195 -7836 -1185 -7676
rect -1133 -7836 -1123 -7676
rect -1084 -7824 -1078 -7596
rect -1044 -7824 -1038 -7596
rect -986 -7676 -980 -7448
rect -946 -7676 -940 -7448
rect -901 -7596 -891 -7436
rect -839 -7596 -829 -7436
rect -790 -7448 -744 -7436
rect -1084 -7836 -1038 -7824
rect -999 -7836 -989 -7676
rect -937 -7836 -927 -7676
rect -888 -7824 -882 -7596
rect -848 -7824 -842 -7596
rect -790 -7676 -784 -7448
rect -750 -7676 -744 -7448
rect -705 -7596 -695 -7436
rect -643 -7596 -633 -7436
rect -594 -7448 -548 -7436
rect -888 -7836 -842 -7824
rect -803 -7836 -793 -7676
rect -741 -7836 -731 -7676
rect -692 -7824 -686 -7596
rect -652 -7824 -646 -7596
rect -594 -7676 -588 -7448
rect -554 -7676 -548 -7448
rect -509 -7596 -499 -7436
rect -447 -7596 -437 -7436
rect -398 -7448 -352 -7436
rect -692 -7836 -646 -7824
rect -607 -7836 -597 -7676
rect -545 -7836 -535 -7676
rect -496 -7824 -490 -7596
rect -456 -7824 -450 -7596
rect -398 -7676 -392 -7448
rect -358 -7676 -352 -7448
rect -313 -7596 -303 -7436
rect -251 -7596 -241 -7436
rect -202 -7448 -156 -7436
rect -496 -7836 -450 -7824
rect -411 -7836 -401 -7676
rect -349 -7836 -339 -7676
rect -300 -7824 -294 -7596
rect -260 -7824 -254 -7596
rect -202 -7676 -196 -7448
rect -162 -7676 -156 -7448
rect -117 -7596 -107 -7436
rect -55 -7596 -45 -7436
rect -6 -7448 40 -7436
rect -300 -7836 -254 -7824
rect -215 -7836 -205 -7676
rect -153 -7836 -143 -7676
rect -104 -7824 -98 -7596
rect -64 -7824 -58 -7596
rect -6 -7676 0 -7448
rect 34 -7676 40 -7448
rect 79 -7596 89 -7436
rect 141 -7596 151 -7436
rect 190 -7448 236 -7436
rect -104 -7836 -58 -7824
rect -19 -7836 -9 -7676
rect 43 -7836 53 -7676
rect 92 -7824 98 -7596
rect 132 -7824 138 -7596
rect 190 -7676 196 -7448
rect 230 -7676 236 -7448
rect 275 -7596 285 -7436
rect 337 -7596 347 -7436
rect 386 -7448 432 -7436
rect 92 -7836 138 -7824
rect 177 -7836 187 -7676
rect 239 -7836 249 -7676
rect 288 -7824 294 -7596
rect 328 -7824 334 -7596
rect 386 -7676 392 -7448
rect 426 -7676 432 -7448
rect 471 -7596 481 -7436
rect 533 -7596 543 -7436
rect 582 -7448 628 -7436
rect 288 -7836 334 -7824
rect 373 -7836 383 -7676
rect 435 -7836 445 -7676
rect 484 -7824 490 -7596
rect 524 -7824 530 -7596
rect 582 -7676 588 -7448
rect 622 -7676 628 -7448
rect 667 -7596 677 -7436
rect 729 -7596 739 -7436
rect 778 -7448 824 -7436
rect 484 -7836 530 -7824
rect 569 -7836 579 -7676
rect 631 -7836 641 -7676
rect 680 -7824 686 -7596
rect 720 -7824 726 -7596
rect 778 -7676 784 -7448
rect 818 -7676 824 -7448
rect 863 -7596 873 -7436
rect 925 -7596 935 -7436
rect 974 -7448 1020 -7436
rect 680 -7836 726 -7824
rect 765 -7836 775 -7676
rect 827 -7836 837 -7676
rect 876 -7824 882 -7596
rect 916 -7824 922 -7596
rect 974 -7676 980 -7448
rect 1014 -7676 1020 -7448
rect 1059 -7596 1069 -7436
rect 1121 -7596 1131 -7436
rect 1170 -7448 1216 -7436
rect 876 -7836 922 -7824
rect 961 -7836 971 -7676
rect 1023 -7836 1033 -7676
rect 1072 -7824 1078 -7596
rect 1112 -7824 1118 -7596
rect 1170 -7676 1176 -7448
rect 1210 -7676 1216 -7448
rect 1255 -7596 1265 -7436
rect 1317 -7596 1327 -7436
rect 1072 -7836 1118 -7824
rect 1157 -7836 1167 -7676
rect 1219 -7836 1229 -7676
rect 1268 -7824 1274 -7596
rect 1308 -7824 1314 -7596
rect 1268 -7836 1314 -7824
rect -1144 -7870 1274 -7864
rect 1404 -7870 1544 -7400
rect 2344 -7360 2434 -6890
rect 2517 -6892 2533 -6890
rect 2567 -6892 2631 -6858
rect 2665 -6892 2729 -6858
rect 2763 -6892 2827 -6858
rect 2861 -6892 2925 -6858
rect 2959 -6892 3023 -6858
rect 3057 -6892 3121 -6858
rect 3155 -6892 3219 -6858
rect 3253 -6892 3317 -6858
rect 3351 -6892 3415 -6858
rect 3449 -6892 3513 -6858
rect 3547 -6892 3611 -6858
rect 3645 -6892 3709 -6858
rect 3743 -6892 3807 -6858
rect 3841 -6892 3905 -6858
rect 3939 -6892 3955 -6858
rect 2517 -6898 3955 -6892
rect 2478 -6942 2524 -6930
rect 2478 -7170 2484 -6942
rect 2518 -7170 2524 -6942
rect 2563 -7090 2573 -6930
rect 2625 -7090 2635 -6930
rect 2674 -6942 2720 -6930
rect 2465 -7330 2475 -7170
rect 2527 -7330 2537 -7170
rect 2576 -7318 2582 -7090
rect 2616 -7318 2622 -7090
rect 2674 -7170 2680 -6942
rect 2714 -7170 2720 -6942
rect 2759 -7090 2769 -6930
rect 2821 -7090 2831 -6930
rect 2870 -6942 2916 -6930
rect 2576 -7330 2622 -7318
rect 2661 -7330 2671 -7170
rect 2723 -7330 2733 -7170
rect 2772 -7318 2778 -7090
rect 2812 -7318 2818 -7090
rect 2870 -7170 2876 -6942
rect 2910 -7170 2916 -6942
rect 2955 -7090 2965 -6930
rect 3017 -7090 3027 -6930
rect 3066 -6942 3112 -6930
rect 2772 -7330 2818 -7318
rect 2857 -7330 2867 -7170
rect 2919 -7330 2929 -7170
rect 2968 -7318 2974 -7090
rect 3008 -7318 3014 -7090
rect 3066 -7170 3072 -6942
rect 3106 -7170 3112 -6942
rect 3151 -7090 3161 -6930
rect 3213 -7090 3223 -6930
rect 3262 -6942 3308 -6930
rect 2968 -7330 3014 -7318
rect 3053 -7330 3063 -7170
rect 3115 -7330 3125 -7170
rect 3164 -7318 3170 -7090
rect 3204 -7318 3210 -7090
rect 3262 -7170 3268 -6942
rect 3302 -7170 3308 -6942
rect 3347 -7090 3357 -6930
rect 3409 -7090 3419 -6930
rect 3458 -6942 3504 -6930
rect 3164 -7330 3210 -7318
rect 3249 -7330 3259 -7170
rect 3311 -7330 3321 -7170
rect 3360 -7318 3366 -7090
rect 3400 -7318 3406 -7090
rect 3458 -7170 3464 -6942
rect 3498 -7170 3504 -6942
rect 3543 -7090 3553 -6930
rect 3605 -7090 3615 -6930
rect 3654 -6942 3700 -6930
rect 3360 -7330 3406 -7318
rect 3445 -7330 3455 -7170
rect 3507 -7330 3517 -7170
rect 3556 -7318 3562 -7090
rect 3596 -7318 3602 -7090
rect 3654 -7170 3660 -6942
rect 3694 -7170 3700 -6942
rect 3739 -7090 3749 -6930
rect 3801 -7090 3811 -6930
rect 3850 -6942 3896 -6930
rect 3556 -7330 3602 -7318
rect 3641 -7330 3651 -7170
rect 3703 -7330 3713 -7170
rect 3752 -7318 3758 -7090
rect 3792 -7318 3798 -7090
rect 3850 -7170 3856 -6942
rect 3890 -7170 3896 -6942
rect 3935 -7090 3945 -6930
rect 3997 -7090 4007 -6930
rect 4044 -6940 4054 -6730
rect 4174 -6940 4184 -6730
rect 4048 -6952 4180 -6940
rect 3752 -7330 3798 -7318
rect 3837 -7330 3847 -7170
rect 3899 -7330 3909 -7170
rect 3948 -7318 3954 -7090
rect 3988 -7318 3994 -7090
rect 3948 -7330 3994 -7318
rect 2344 -7362 2524 -7360
rect 2344 -7368 3955 -7362
rect 2344 -7402 2533 -7368
rect 2567 -7402 2631 -7368
rect 2665 -7402 2729 -7368
rect 2763 -7402 2827 -7368
rect 2861 -7402 2925 -7368
rect 2959 -7402 3023 -7368
rect 3057 -7402 3121 -7368
rect 3155 -7402 3219 -7368
rect 3253 -7402 3317 -7368
rect 3351 -7402 3415 -7368
rect 3449 -7402 3513 -7368
rect 3547 -7402 3611 -7368
rect 3645 -7402 3709 -7368
rect 3743 -7402 3807 -7368
rect 3841 -7402 3905 -7368
rect 3939 -7402 3955 -7368
rect 2344 -7418 3955 -7402
rect 2344 -7420 2524 -7418
rect -1386 -7874 1544 -7870
rect -1386 -7908 -1128 -7874
rect -1094 -7908 -1029 -7874
rect -995 -7908 -932 -7874
rect -898 -7908 -833 -7874
rect -799 -7908 -736 -7874
rect -702 -7908 -637 -7874
rect -603 -7908 -540 -7874
rect -506 -7908 -441 -7874
rect -407 -7908 -344 -7874
rect -310 -7908 -245 -7874
rect -211 -7908 -148 -7874
rect -114 -7908 -49 -7874
rect -15 -7908 48 -7874
rect 82 -7908 147 -7874
rect 181 -7908 244 -7874
rect 278 -7908 343 -7874
rect 377 -7908 440 -7874
rect 474 -7908 539 -7874
rect 573 -7908 636 -7874
rect 670 -7908 735 -7874
rect 769 -7908 832 -7874
rect 866 -7908 931 -7874
rect 965 -7908 1028 -7874
rect 1062 -7908 1127 -7874
rect 1161 -7908 1224 -7874
rect 1258 -7908 1544 -7874
rect -1386 -7982 1544 -7908
rect -1386 -8016 -1127 -7982
rect -1093 -8016 -1029 -7982
rect -995 -8016 -931 -7982
rect -897 -8016 -833 -7982
rect -799 -8016 -735 -7982
rect -701 -8016 -637 -7982
rect -603 -8016 -539 -7982
rect -505 -8016 -441 -7982
rect -407 -8016 -343 -7982
rect -309 -8016 -245 -7982
rect -211 -8016 -147 -7982
rect -113 -8016 -49 -7982
rect -15 -8016 49 -7982
rect 83 -8016 147 -7982
rect 181 -8016 245 -7982
rect 279 -8016 343 -7982
rect 377 -8016 441 -7982
rect 475 -8016 539 -7982
rect 573 -8016 637 -7982
rect 671 -8016 735 -7982
rect 769 -8016 833 -7982
rect 867 -8016 931 -7982
rect 965 -8016 1029 -7982
rect 1063 -8016 1127 -7982
rect 1161 -8016 1225 -7982
rect 1259 -8016 1544 -7982
rect 4470 -7990 4620 -2350
rect -1386 -8020 1544 -8016
rect -1386 -8490 -1236 -8020
rect -1143 -8026 1275 -8020
rect -1195 -8214 -1185 -8054
rect -1133 -8214 -1123 -8054
rect -1084 -8066 -1038 -8054
rect -1182 -8442 -1176 -8214
rect -1142 -8442 -1136 -8214
rect -1084 -8294 -1078 -8066
rect -1044 -8294 -1038 -8066
rect -999 -8214 -989 -8054
rect -937 -8214 -927 -8054
rect -888 -8066 -842 -8054
rect -1182 -8454 -1136 -8442
rect -1097 -8454 -1087 -8294
rect -1035 -8454 -1025 -8294
rect -986 -8442 -980 -8214
rect -946 -8442 -940 -8214
rect -888 -8294 -882 -8066
rect -848 -8294 -842 -8066
rect -803 -8214 -793 -8054
rect -741 -8214 -731 -8054
rect -692 -8066 -646 -8054
rect -986 -8454 -940 -8442
rect -901 -8454 -891 -8294
rect -839 -8454 -829 -8294
rect -790 -8442 -784 -8214
rect -750 -8442 -744 -8214
rect -692 -8294 -686 -8066
rect -652 -8294 -646 -8066
rect -607 -8214 -597 -8054
rect -545 -8214 -535 -8054
rect -496 -8066 -450 -8054
rect -790 -8454 -744 -8442
rect -705 -8454 -695 -8294
rect -643 -8454 -633 -8294
rect -594 -8442 -588 -8214
rect -554 -8442 -548 -8214
rect -496 -8294 -490 -8066
rect -456 -8294 -450 -8066
rect -411 -8214 -401 -8054
rect -349 -8214 -339 -8054
rect -300 -8066 -254 -8054
rect -594 -8454 -548 -8442
rect -509 -8454 -499 -8294
rect -447 -8454 -437 -8294
rect -398 -8442 -392 -8214
rect -358 -8442 -352 -8214
rect -300 -8294 -294 -8066
rect -260 -8294 -254 -8066
rect -215 -8214 -205 -8054
rect -153 -8214 -143 -8054
rect -104 -8066 -58 -8054
rect -398 -8454 -352 -8442
rect -313 -8454 -303 -8294
rect -251 -8454 -241 -8294
rect -202 -8442 -196 -8214
rect -162 -8442 -156 -8214
rect -104 -8294 -98 -8066
rect -64 -8294 -58 -8066
rect -19 -8214 -9 -8054
rect 43 -8214 53 -8054
rect 92 -8066 138 -8054
rect -202 -8454 -156 -8442
rect -117 -8454 -107 -8294
rect -55 -8454 -45 -8294
rect -6 -8442 0 -8214
rect 34 -8442 40 -8214
rect 92 -8294 98 -8066
rect 132 -8294 138 -8066
rect 177 -8214 187 -8054
rect 239 -8214 249 -8054
rect 288 -8066 334 -8054
rect -6 -8454 40 -8442
rect 79 -8454 89 -8294
rect 141 -8454 151 -8294
rect 190 -8442 196 -8214
rect 230 -8442 236 -8214
rect 288 -8294 294 -8066
rect 328 -8294 334 -8066
rect 373 -8214 383 -8054
rect 435 -8214 445 -8054
rect 484 -8066 530 -8054
rect 190 -8454 236 -8442
rect 275 -8454 285 -8294
rect 337 -8454 347 -8294
rect 386 -8442 392 -8214
rect 426 -8442 432 -8214
rect 484 -8294 490 -8066
rect 524 -8294 530 -8066
rect 569 -8214 579 -8054
rect 631 -8214 641 -8054
rect 680 -8066 726 -8054
rect 386 -8454 432 -8442
rect 471 -8454 481 -8294
rect 533 -8454 543 -8294
rect 582 -8442 588 -8214
rect 622 -8442 628 -8214
rect 680 -8294 686 -8066
rect 720 -8294 726 -8066
rect 765 -8214 775 -8054
rect 827 -8214 837 -8054
rect 876 -8066 922 -8054
rect 582 -8454 628 -8442
rect 667 -8454 677 -8294
rect 729 -8454 739 -8294
rect 778 -8442 784 -8214
rect 818 -8442 824 -8214
rect 876 -8294 882 -8066
rect 916 -8294 922 -8066
rect 961 -8214 971 -8054
rect 1023 -8214 1033 -8054
rect 1072 -8066 1118 -8054
rect 778 -8454 824 -8442
rect 863 -8454 873 -8294
rect 925 -8454 935 -8294
rect 974 -8442 980 -8214
rect 1014 -8442 1020 -8214
rect 1072 -8294 1078 -8066
rect 1112 -8294 1118 -8066
rect 1157 -8214 1167 -8054
rect 1219 -8214 1229 -8054
rect 1268 -8066 1314 -8054
rect 974 -8454 1020 -8442
rect 1059 -8454 1069 -8294
rect 1121 -8454 1131 -8294
rect 1170 -8442 1176 -8214
rect 1210 -8442 1216 -8214
rect 1268 -8294 1274 -8066
rect 1308 -8294 1314 -8066
rect 1170 -8454 1216 -8442
rect 1255 -8454 1265 -8294
rect 1317 -8454 1327 -8294
rect 1404 -8480 1544 -8020
rect 1644 -8018 2850 -7990
rect 1644 -8052 1662 -8018
rect 1696 -8052 1758 -8018
rect 1792 -8052 1854 -8018
rect 1888 -8052 1950 -8018
rect 1984 -8052 2046 -8018
rect 2080 -8052 2142 -8018
rect 2176 -8052 2238 -8018
rect 2272 -8052 2334 -8018
rect 2368 -8052 2430 -8018
rect 2464 -8052 2526 -8018
rect 2560 -8052 2622 -8018
rect 2656 -8052 2718 -8018
rect 2752 -8052 2850 -8018
rect 1644 -8060 2850 -8052
rect 1608 -8102 1654 -8090
rect 1608 -8330 1614 -8102
rect 1648 -8330 1654 -8102
rect 1691 -8250 1701 -8090
rect 1753 -8250 1763 -8090
rect 1800 -8102 1846 -8090
rect -1143 -8490 1275 -8482
rect 1384 -8490 1544 -8480
rect 1595 -8490 1605 -8330
rect 1657 -8490 1667 -8330
rect 1704 -8478 1710 -8250
rect 1744 -8478 1750 -8250
rect 1800 -8330 1806 -8102
rect 1840 -8330 1846 -8102
rect 1883 -8250 1893 -8090
rect 1945 -8250 1955 -8090
rect 1992 -8102 2038 -8090
rect 1704 -8490 1750 -8478
rect 1787 -8490 1797 -8330
rect 1849 -8490 1859 -8330
rect 1896 -8478 1902 -8250
rect 1936 -8478 1942 -8250
rect 1992 -8330 1998 -8102
rect 2032 -8330 2038 -8102
rect 2075 -8250 2085 -8090
rect 2137 -8250 2147 -8090
rect 2184 -8102 2230 -8090
rect 1896 -8490 1942 -8478
rect 1979 -8490 1989 -8330
rect 2041 -8490 2051 -8330
rect 2088 -8478 2094 -8250
rect 2128 -8478 2134 -8250
rect 2184 -8330 2190 -8102
rect 2224 -8330 2230 -8102
rect 2267 -8250 2277 -8090
rect 2329 -8250 2339 -8090
rect 2376 -8102 2422 -8090
rect 2088 -8490 2134 -8478
rect 2171 -8490 2181 -8330
rect 2233 -8490 2243 -8330
rect 2280 -8478 2286 -8250
rect 2320 -8478 2326 -8250
rect 2376 -8330 2382 -8102
rect 2416 -8330 2422 -8102
rect 2459 -8250 2469 -8090
rect 2521 -8250 2531 -8090
rect 2568 -8102 2614 -8090
rect 2280 -8490 2326 -8478
rect 2363 -8490 2373 -8330
rect 2425 -8490 2435 -8330
rect 2472 -8478 2478 -8250
rect 2512 -8478 2518 -8250
rect 2568 -8330 2574 -8102
rect 2608 -8330 2614 -8102
rect 2651 -8250 2661 -8090
rect 2713 -8250 2723 -8090
rect 2760 -8102 2806 -8090
rect 2472 -8490 2518 -8478
rect 2555 -8490 2565 -8330
rect 2617 -8490 2627 -8330
rect 2664 -8478 2670 -8250
rect 2704 -8478 2710 -8250
rect 2760 -8330 2766 -8102
rect 2800 -8330 2806 -8102
rect 2840 -8140 2850 -8060
rect 3020 -8140 3030 -7990
rect 3540 -8018 4860 -7990
rect 3540 -8052 3558 -8018
rect 3592 -8052 3654 -8018
rect 3688 -8052 3750 -8018
rect 3784 -8052 3846 -8018
rect 3880 -8052 3942 -8018
rect 3976 -8052 4038 -8018
rect 4072 -8052 4134 -8018
rect 4168 -8052 4230 -8018
rect 4264 -8052 4326 -8018
rect 4360 -8052 4422 -8018
rect 4456 -8052 4518 -8018
rect 4552 -8052 4614 -8018
rect 4648 -8052 4860 -8018
rect 3540 -8060 4860 -8052
rect 3600 -8090 3650 -8060
rect 3790 -8090 3840 -8060
rect 3980 -8090 4030 -8060
rect 4170 -8090 4220 -8060
rect 4370 -8090 4420 -8060
rect 4560 -8090 4610 -8060
rect 3504 -8102 3550 -8090
rect 2664 -8490 2710 -8478
rect 2747 -8490 2757 -8330
rect 2809 -8490 2819 -8330
rect -1386 -8492 1544 -8490
rect -1386 -8526 -1127 -8492
rect -1093 -8526 -1029 -8492
rect -995 -8526 -931 -8492
rect -897 -8526 -833 -8492
rect -799 -8526 -735 -8492
rect -701 -8526 -637 -8492
rect -603 -8526 -539 -8492
rect -505 -8526 -441 -8492
rect -407 -8526 -343 -8492
rect -309 -8526 -245 -8492
rect -211 -8526 -147 -8492
rect -113 -8526 -49 -8492
rect -15 -8526 49 -8492
rect 83 -8526 147 -8492
rect 181 -8526 245 -8492
rect 279 -8526 343 -8492
rect 377 -8526 441 -8492
rect 475 -8526 539 -8492
rect 573 -8526 637 -8492
rect 671 -8526 735 -8492
rect 769 -8526 833 -8492
rect 867 -8526 931 -8492
rect 965 -8526 1029 -8492
rect 1063 -8526 1127 -8492
rect 1161 -8526 1225 -8492
rect 1259 -8526 1544 -8492
rect 2854 -8520 2964 -8140
rect 3504 -8330 3510 -8102
rect 3544 -8330 3550 -8102
rect 3587 -8250 3597 -8090
rect 3649 -8250 3659 -8090
rect 3696 -8102 3742 -8090
rect 3491 -8490 3501 -8330
rect 3553 -8490 3563 -8330
rect 3600 -8478 3606 -8250
rect 3640 -8478 3646 -8250
rect 3696 -8330 3702 -8102
rect 3736 -8330 3742 -8102
rect 3779 -8250 3789 -8090
rect 3841 -8250 3851 -8090
rect 3888 -8102 3934 -8090
rect 3600 -8490 3646 -8478
rect 3683 -8490 3693 -8330
rect 3745 -8490 3755 -8330
rect 3792 -8478 3798 -8250
rect 3832 -8478 3838 -8250
rect 3888 -8330 3894 -8102
rect 3928 -8330 3934 -8102
rect 3971 -8250 3981 -8090
rect 4033 -8250 4043 -8090
rect 4080 -8102 4126 -8090
rect 3792 -8490 3838 -8478
rect 3875 -8490 3885 -8330
rect 3937 -8490 3947 -8330
rect 3984 -8478 3990 -8250
rect 4024 -8478 4030 -8250
rect 4080 -8330 4086 -8102
rect 4120 -8330 4126 -8102
rect 4163 -8250 4173 -8090
rect 4225 -8250 4235 -8090
rect 4272 -8102 4318 -8090
rect 3984 -8490 4030 -8478
rect 4067 -8490 4077 -8330
rect 4129 -8490 4139 -8330
rect 4176 -8478 4182 -8250
rect 4216 -8478 4222 -8250
rect 4272 -8330 4278 -8102
rect 4312 -8330 4318 -8102
rect 4355 -8250 4365 -8090
rect 4417 -8250 4427 -8090
rect 4464 -8102 4510 -8090
rect 4176 -8490 4222 -8478
rect 4259 -8490 4269 -8330
rect 4321 -8490 4331 -8330
rect 4368 -8478 4374 -8250
rect 4408 -8478 4414 -8250
rect 4464 -8330 4470 -8102
rect 4504 -8330 4510 -8102
rect 4547 -8250 4557 -8090
rect 4609 -8250 4619 -8090
rect 4656 -8102 4702 -8090
rect 4368 -8490 4414 -8478
rect 4451 -8490 4461 -8330
rect 4513 -8490 4523 -8330
rect 4560 -8478 4566 -8250
rect 4600 -8478 4606 -8250
rect 4656 -8330 4662 -8102
rect 4696 -8330 4702 -8102
rect 4560 -8490 4606 -8478
rect 4643 -8490 4653 -8330
rect 4705 -8490 4715 -8330
rect 4750 -8520 4860 -8060
rect -1386 -8540 1544 -8526
rect 1644 -8528 2964 -8520
rect -1143 -8542 1275 -8540
rect 1644 -8562 1662 -8528
rect 1696 -8562 1758 -8528
rect 1792 -8562 1854 -8528
rect 1888 -8562 1950 -8528
rect 1984 -8562 2046 -8528
rect 2080 -8562 2142 -8528
rect 2176 -8562 2238 -8528
rect 2272 -8562 2334 -8528
rect 2368 -8562 2430 -8528
rect 2464 -8562 2526 -8528
rect 2560 -8562 2622 -8528
rect 2656 -8562 2718 -8528
rect 2752 -8562 2964 -8528
rect 1644 -8590 2964 -8562
rect 3540 -8528 4860 -8520
rect 3540 -8562 3558 -8528
rect 3592 -8562 3654 -8528
rect 3688 -8562 3750 -8528
rect 3784 -8562 3846 -8528
rect 3880 -8562 3942 -8528
rect 3976 -8562 4038 -8528
rect 4072 -8562 4134 -8528
rect 4168 -8562 4230 -8528
rect 4264 -8562 4326 -8528
rect 4360 -8562 4422 -8528
rect 4456 -8562 4518 -8528
rect 4552 -8562 4614 -8528
rect 4648 -8562 4860 -8528
rect 3540 -8590 4860 -8562
rect -1390 -8850 -1380 -8760
rect -1270 -8767 -1196 -8760
rect -1270 -8784 1247 -8767
rect -1270 -8818 -1148 -8784
rect -1114 -8818 -956 -8784
rect -922 -8818 -764 -8784
rect -730 -8818 -572 -8784
rect -538 -8818 -380 -8784
rect -346 -8818 -188 -8784
rect -154 -8818 4 -8784
rect 38 -8818 196 -8784
rect 230 -8818 388 -8784
rect 422 -8818 580 -8784
rect 614 -8818 772 -8784
rect 806 -8818 964 -8784
rect 998 -8818 1156 -8784
rect 1190 -8818 1247 -8784
rect 2834 -8800 2964 -8590
rect 4730 -8800 4860 -8590
rect -1270 -8820 1247 -8818
rect -1270 -8850 -1246 -8820
rect -1203 -8827 1247 -8820
rect -1346 -9290 -1246 -8850
rect 1654 -8838 5480 -8800
rect -1202 -8868 -1156 -8856
rect -1202 -9096 -1196 -8868
rect -1162 -9096 -1156 -8868
rect -1119 -9016 -1109 -8856
rect -1057 -9016 -1047 -8856
rect -1010 -8868 -964 -8856
rect -1215 -9256 -1205 -9096
rect -1153 -9256 -1143 -9096
rect -1106 -9244 -1100 -9016
rect -1066 -9244 -1060 -9016
rect -1010 -9096 -1004 -8868
rect -970 -9096 -964 -8868
rect -927 -9016 -917 -8856
rect -865 -9016 -855 -8856
rect -818 -8868 -772 -8856
rect -1106 -9256 -1060 -9244
rect -1023 -9256 -1013 -9096
rect -961 -9256 -951 -9096
rect -914 -9244 -908 -9016
rect -874 -9244 -868 -9016
rect -818 -9096 -812 -8868
rect -778 -9096 -772 -8868
rect -735 -9016 -725 -8856
rect -673 -9016 -663 -8856
rect -626 -8868 -580 -8856
rect -914 -9256 -868 -9244
rect -831 -9256 -821 -9096
rect -769 -9256 -759 -9096
rect -722 -9244 -716 -9016
rect -682 -9244 -676 -9016
rect -626 -9096 -620 -8868
rect -586 -9096 -580 -8868
rect -543 -9016 -533 -8856
rect -481 -9016 -471 -8856
rect -434 -8868 -388 -8856
rect -722 -9256 -676 -9244
rect -639 -9256 -629 -9096
rect -577 -9256 -567 -9096
rect -530 -9244 -524 -9016
rect -490 -9244 -484 -9016
rect -434 -9096 -428 -8868
rect -394 -9096 -388 -8868
rect -351 -9016 -341 -8856
rect -289 -9016 -279 -8856
rect -242 -8868 -196 -8856
rect -530 -9256 -484 -9244
rect -447 -9256 -437 -9096
rect -385 -9256 -375 -9096
rect -338 -9244 -332 -9016
rect -298 -9244 -292 -9016
rect -242 -9096 -236 -8868
rect -202 -9096 -196 -8868
rect -159 -9016 -149 -8856
rect -97 -9016 -87 -8856
rect -50 -8868 -4 -8856
rect -338 -9256 -292 -9244
rect -255 -9256 -245 -9096
rect -193 -9256 -183 -9096
rect -146 -9244 -140 -9016
rect -106 -9244 -100 -9016
rect -50 -9096 -44 -8868
rect -10 -9096 -4 -8868
rect 33 -9016 43 -8856
rect 95 -9016 105 -8856
rect 142 -8868 188 -8856
rect -146 -9256 -100 -9244
rect -63 -9256 -53 -9096
rect -1 -9256 9 -9096
rect 46 -9244 52 -9016
rect 86 -9244 92 -9016
rect 142 -9096 148 -8868
rect 182 -9096 188 -8868
rect 225 -9016 235 -8856
rect 287 -9016 297 -8856
rect 334 -8868 380 -8856
rect 46 -9256 92 -9244
rect 129 -9256 139 -9096
rect 191 -9256 201 -9096
rect 238 -9244 244 -9016
rect 278 -9244 284 -9016
rect 334 -9096 340 -8868
rect 374 -9096 380 -8868
rect 417 -9016 427 -8856
rect 479 -9016 489 -8856
rect 526 -8868 572 -8856
rect 238 -9256 284 -9244
rect 321 -9256 331 -9096
rect 383 -9256 393 -9096
rect 430 -9244 436 -9016
rect 470 -9244 476 -9016
rect 526 -9096 532 -8868
rect 566 -9096 572 -8868
rect 609 -9016 619 -8856
rect 671 -9016 681 -8856
rect 718 -8868 764 -8856
rect 430 -9256 476 -9244
rect 513 -9256 523 -9096
rect 575 -9256 585 -9096
rect 622 -9244 628 -9016
rect 662 -9244 668 -9016
rect 718 -9096 724 -8868
rect 758 -9096 764 -8868
rect 801 -9016 811 -8856
rect 863 -9016 873 -8856
rect 910 -8868 956 -8856
rect 622 -9256 668 -9244
rect 705 -9256 715 -9096
rect 767 -9256 777 -9096
rect 814 -9244 820 -9016
rect 854 -9244 860 -9016
rect 910 -9096 916 -8868
rect 950 -9096 956 -8868
rect 993 -9016 1003 -8856
rect 1055 -9016 1065 -8856
rect 1102 -8868 1148 -8856
rect 814 -9256 860 -9244
rect 897 -9256 907 -9096
rect 959 -9256 969 -9096
rect 1006 -9244 1012 -9016
rect 1046 -9244 1052 -9016
rect 1102 -9096 1108 -8868
rect 1142 -9096 1148 -8868
rect 1185 -9016 1195 -8856
rect 1247 -9016 1257 -8856
rect 1654 -8872 1676 -8838
rect 1844 -8872 1934 -8838
rect 2102 -8872 2192 -8838
rect 2360 -8872 2450 -8838
rect 2618 -8872 2708 -8838
rect 2876 -8872 2966 -8838
rect 3134 -8872 3572 -8838
rect 3740 -8872 3830 -8838
rect 3998 -8872 4088 -8838
rect 4256 -8872 4346 -8838
rect 4514 -8872 4604 -8838
rect 4772 -8872 4862 -8838
rect 5030 -8872 5480 -8838
rect 1654 -8880 5480 -8872
rect 5590 -8838 6130 -8810
rect 5590 -8872 5604 -8838
rect 5638 -8872 5796 -8838
rect 5830 -8872 6130 -8838
rect 5590 -8880 6130 -8872
rect 1608 -8922 1654 -8910
rect 1006 -9256 1052 -9244
rect 1089 -9256 1099 -9096
rect 1151 -9256 1161 -9096
rect 1198 -9244 1204 -9016
rect 1238 -9244 1244 -9016
rect 1338 -9140 1480 -9128
rect 1198 -9256 1244 -9244
rect -1203 -9290 1247 -9287
rect -1346 -9294 1247 -9290
rect -1346 -9328 -1052 -9294
rect -1018 -9328 -860 -9294
rect -826 -9328 -668 -9294
rect -634 -9328 -476 -9294
rect -442 -9328 -284 -9294
rect -250 -9328 -92 -9294
rect -58 -9328 100 -9294
rect 134 -9328 292 -9294
rect 326 -9328 484 -9294
rect 518 -9328 676 -9294
rect 710 -9328 868 -9294
rect 902 -9328 1060 -9294
rect 1094 -9328 1247 -9294
rect 1334 -9320 1344 -9140
rect 1474 -9320 1484 -9140
rect 1608 -9150 1614 -8922
rect 1648 -9150 1654 -8922
rect 1853 -9070 1863 -8910
rect 1915 -9070 1925 -8910
rect 2124 -8922 2170 -8910
rect 1595 -9310 1605 -9150
rect 1657 -9310 1667 -9150
rect 1866 -9298 1872 -9070
rect 1906 -9298 1912 -9070
rect 2124 -9150 2130 -8922
rect 2164 -9150 2170 -8922
rect 2369 -9070 2379 -8910
rect 2431 -9070 2441 -8910
rect 2640 -8922 2686 -8910
rect 1866 -9310 1912 -9298
rect 2111 -9310 2121 -9150
rect 2173 -9310 2183 -9150
rect 2382 -9298 2388 -9070
rect 2422 -9298 2428 -9070
rect 2640 -9150 2646 -8922
rect 2680 -9150 2686 -8922
rect 2885 -9070 2895 -8910
rect 2947 -9070 2954 -8910
rect 2382 -9310 2428 -9298
rect 2627 -9310 2637 -9150
rect 2689 -9310 2699 -9150
rect 2898 -9298 2904 -9070
rect 2938 -9298 2944 -9070
rect 2898 -9310 2944 -9298
rect -1346 -9402 1247 -9328
rect 1338 -9332 1480 -9320
rect 3004 -9340 3094 -8880
rect 3156 -8922 3202 -8910
rect 3156 -9150 3162 -8922
rect 3196 -9150 3202 -8922
rect 3504 -8922 3550 -8910
rect 3504 -9150 3510 -8922
rect 3544 -9150 3550 -8922
rect 3749 -9070 3759 -8910
rect 3811 -9070 3821 -8910
rect 4020 -8922 4066 -8910
rect 3143 -9310 3153 -9150
rect 3205 -9310 3215 -9150
rect 3491 -9310 3501 -9150
rect 3553 -9310 3563 -9150
rect 3762 -9298 3768 -9070
rect 3802 -9298 3808 -9070
rect 4020 -9150 4026 -8922
rect 4060 -9150 4066 -8922
rect 4265 -9070 4275 -8910
rect 4327 -9070 4337 -8910
rect 4536 -8922 4582 -8910
rect 3762 -9310 3808 -9298
rect 4007 -9310 4017 -9150
rect 4069 -9310 4079 -9150
rect 4278 -9298 4284 -9070
rect 4318 -9298 4324 -9070
rect 4536 -9150 4542 -8922
rect 4576 -9150 4582 -8922
rect 4781 -9070 4791 -8910
rect 4843 -9070 4850 -8910
rect 4278 -9310 4324 -9298
rect 4523 -9310 4533 -9150
rect 4585 -9310 4595 -9150
rect 4794 -9298 4800 -9070
rect 4834 -9298 4840 -9070
rect 4794 -9310 4840 -9298
rect 4900 -9340 4990 -8880
rect 5390 -8910 5480 -8880
rect 5052 -8922 5098 -8910
rect 5052 -9150 5058 -8922
rect 5092 -9150 5098 -8922
rect 5390 -9090 5440 -8910
rect 5500 -9090 5510 -8910
rect 5550 -8922 5596 -8910
rect 5039 -9310 5049 -9150
rect 5101 -9310 5111 -9150
rect 5454 -9298 5460 -9090
rect 5494 -9298 5500 -9090
rect 5550 -9150 5556 -8922
rect 5590 -9150 5596 -8922
rect 5630 -9090 5640 -8910
rect 5700 -9090 5710 -8910
rect 5742 -8922 5788 -8910
rect 5454 -9310 5500 -9298
rect 5530 -9310 5540 -9150
rect 5600 -9310 5610 -9150
rect 5646 -9298 5652 -9090
rect 5686 -9298 5692 -9090
rect 5742 -9150 5748 -8922
rect 5782 -9150 5788 -8922
rect 5820 -9090 5830 -8910
rect 5890 -9090 5900 -8910
rect 5934 -8922 5980 -8910
rect 5646 -9310 5692 -9298
rect 5730 -9310 5740 -9150
rect 5800 -9310 5810 -9150
rect 5838 -9298 5844 -9090
rect 5878 -9298 5884 -9090
rect 5934 -9150 5940 -8922
rect 5974 -9150 5980 -8922
rect 5838 -9310 5884 -9298
rect 5920 -9310 5930 -9150
rect 5990 -9310 6000 -9150
rect 6030 -9300 6130 -8880
rect 6030 -9340 6060 -9300
rect -1346 -9436 -1052 -9402
rect -1018 -9436 -860 -9402
rect -826 -9436 -668 -9402
rect -634 -9436 -476 -9402
rect -442 -9436 -284 -9402
rect -250 -9436 -92 -9402
rect -58 -9436 100 -9402
rect 134 -9436 292 -9402
rect 326 -9436 484 -9402
rect 518 -9436 676 -9402
rect 710 -9436 868 -9402
rect 902 -9436 1060 -9402
rect 1094 -9436 1247 -9402
rect 1594 -9348 5110 -9340
rect 1594 -9382 1676 -9348
rect 1844 -9382 1934 -9348
rect 2102 -9382 2192 -9348
rect 2360 -9382 2450 -9348
rect 2618 -9382 2708 -9348
rect 2876 -9382 2966 -9348
rect 3134 -9382 3572 -9348
rect 3740 -9382 3830 -9348
rect 3998 -9382 4088 -9348
rect 4256 -9382 4346 -9348
rect 4514 -9382 4604 -9348
rect 4772 -9382 4862 -9348
rect 5030 -9382 5110 -9348
rect 1594 -9420 5110 -9382
rect 5480 -9348 6060 -9340
rect 5480 -9382 5508 -9348
rect 5542 -9382 5700 -9348
rect 5734 -9382 5892 -9348
rect 5926 -9382 6060 -9348
rect 5480 -9410 6060 -9382
rect 6130 -9410 6140 -9300
rect -1346 -9437 1247 -9436
rect -1346 -9440 -1196 -9437
rect -1346 -9910 -1246 -9440
rect -1064 -9442 -1006 -9437
rect -872 -9442 -814 -9437
rect -680 -9442 -622 -9437
rect -488 -9442 -430 -9437
rect -296 -9442 -238 -9437
rect -104 -9442 -46 -9437
rect 88 -9442 146 -9437
rect 280 -9442 338 -9437
rect 472 -9442 530 -9437
rect 664 -9442 722 -9437
rect 856 -9442 914 -9437
rect 1048 -9442 1106 -9437
rect -1215 -9634 -1205 -9474
rect -1153 -9634 -1143 -9474
rect -1106 -9486 -1060 -9474
rect -1202 -9862 -1196 -9634
rect -1162 -9862 -1156 -9634
rect -1106 -9714 -1100 -9486
rect -1066 -9714 -1060 -9486
rect -1023 -9634 -1013 -9474
rect -961 -9634 -951 -9474
rect -914 -9486 -868 -9474
rect -1202 -9874 -1156 -9862
rect -1119 -9874 -1109 -9714
rect -1057 -9874 -1047 -9714
rect -1010 -9862 -1004 -9634
rect -970 -9862 -964 -9634
rect -914 -9714 -908 -9486
rect -874 -9714 -868 -9486
rect -831 -9634 -821 -9474
rect -769 -9634 -759 -9474
rect -722 -9486 -676 -9474
rect -1010 -9874 -964 -9862
rect -927 -9874 -917 -9714
rect -865 -9874 -855 -9714
rect -818 -9862 -812 -9634
rect -778 -9862 -772 -9634
rect -722 -9714 -716 -9486
rect -682 -9714 -676 -9486
rect -639 -9634 -629 -9474
rect -577 -9634 -567 -9474
rect -530 -9486 -484 -9474
rect -818 -9874 -772 -9862
rect -735 -9874 -725 -9714
rect -673 -9874 -663 -9714
rect -626 -9862 -620 -9634
rect -586 -9862 -580 -9634
rect -530 -9714 -524 -9486
rect -490 -9714 -484 -9486
rect -447 -9634 -437 -9474
rect -385 -9634 -375 -9474
rect -338 -9486 -292 -9474
rect -626 -9874 -580 -9862
rect -543 -9874 -533 -9714
rect -481 -9874 -471 -9714
rect -434 -9862 -428 -9634
rect -394 -9862 -388 -9634
rect -338 -9714 -332 -9486
rect -298 -9714 -292 -9486
rect -255 -9634 -245 -9474
rect -193 -9634 -183 -9474
rect -146 -9486 -100 -9474
rect -434 -9874 -388 -9862
rect -351 -9874 -341 -9714
rect -289 -9874 -279 -9714
rect -242 -9862 -236 -9634
rect -202 -9862 -196 -9634
rect -146 -9714 -140 -9486
rect -106 -9714 -100 -9486
rect -63 -9634 -53 -9474
rect -1 -9634 9 -9474
rect 46 -9486 92 -9474
rect -242 -9874 -196 -9862
rect -159 -9874 -149 -9714
rect -97 -9874 -87 -9714
rect -50 -9862 -44 -9634
rect -10 -9862 -4 -9634
rect 46 -9714 52 -9486
rect 86 -9714 92 -9486
rect 129 -9634 139 -9474
rect 191 -9634 201 -9474
rect 238 -9486 284 -9474
rect -50 -9874 -4 -9862
rect 33 -9874 43 -9714
rect 95 -9874 105 -9714
rect 142 -9862 148 -9634
rect 182 -9862 188 -9634
rect 238 -9714 244 -9486
rect 278 -9714 284 -9486
rect 321 -9634 331 -9474
rect 383 -9634 393 -9474
rect 430 -9486 476 -9474
rect 142 -9874 188 -9862
rect 225 -9874 235 -9714
rect 287 -9874 297 -9714
rect 334 -9862 340 -9634
rect 374 -9862 380 -9634
rect 430 -9714 436 -9486
rect 470 -9714 476 -9486
rect 513 -9634 523 -9474
rect 575 -9634 585 -9474
rect 622 -9486 668 -9474
rect 334 -9874 380 -9862
rect 417 -9874 427 -9714
rect 479 -9874 489 -9714
rect 526 -9862 532 -9634
rect 566 -9862 572 -9634
rect 622 -9714 628 -9486
rect 662 -9714 668 -9486
rect 705 -9634 715 -9474
rect 767 -9634 777 -9474
rect 814 -9486 860 -9474
rect 526 -9874 572 -9862
rect 609 -9874 619 -9714
rect 671 -9874 681 -9714
rect 718 -9862 724 -9634
rect 758 -9862 764 -9634
rect 814 -9714 820 -9486
rect 854 -9714 860 -9486
rect 897 -9634 907 -9474
rect 959 -9634 969 -9474
rect 1006 -9486 1052 -9474
rect 718 -9874 764 -9862
rect 801 -9874 811 -9714
rect 863 -9874 873 -9714
rect 910 -9862 916 -9634
rect 950 -9862 956 -9634
rect 1006 -9714 1012 -9486
rect 1046 -9714 1052 -9486
rect 1089 -9634 1099 -9474
rect 1151 -9634 1161 -9474
rect 1198 -9486 1244 -9474
rect 910 -9874 956 -9862
rect 993 -9874 1003 -9714
rect 1055 -9874 1065 -9714
rect 1102 -9862 1108 -9634
rect 1142 -9862 1148 -9634
rect 1198 -9714 1204 -9486
rect 1238 -9714 1244 -9486
rect 1102 -9874 1148 -9862
rect 1185 -9874 1195 -9714
rect 1247 -9874 1257 -9714
rect 1697 -9850 2089 -9844
rect 2617 -9850 3009 -9844
rect 3537 -9850 3929 -9844
rect 4457 -9850 4849 -9844
rect 5377 -9850 5769 -9844
rect 1330 -9884 1709 -9850
rect 2077 -9884 2629 -9850
rect 2997 -9884 3549 -9850
rect 3917 -9884 4469 -9850
rect 4837 -9884 5389 -9850
rect 5757 -9884 6340 -9850
rect 1330 -9890 6340 -9884
rect -1160 -9907 -1102 -9906
rect -968 -9907 -910 -9906
rect -776 -9907 -718 -9906
rect -584 -9907 -526 -9906
rect -392 -9907 -334 -9906
rect -200 -9907 -142 -9906
rect -8 -9907 50 -9906
rect 184 -9907 242 -9906
rect 376 -9907 434 -9906
rect 568 -9907 626 -9906
rect 760 -9907 818 -9906
rect 952 -9907 1010 -9906
rect 1144 -9907 1202 -9906
rect -1203 -9910 1247 -9907
rect 1330 -9910 1380 -9890
rect -1346 -9912 1380 -9910
rect -1346 -9946 -1148 -9912
rect -1114 -9946 -956 -9912
rect -922 -9946 -764 -9912
rect -730 -9946 -572 -9912
rect -538 -9946 -380 -9912
rect -346 -9946 -188 -9912
rect -154 -9946 4 -9912
rect 38 -9946 196 -9912
rect 230 -9946 388 -9912
rect 422 -9946 580 -9912
rect 614 -9946 772 -9912
rect 806 -9946 964 -9912
rect 998 -9946 1156 -9912
rect 1190 -9946 1380 -9912
rect -1346 -10020 1380 -9946
rect -1346 -10054 -1148 -10020
rect -1114 -10054 -956 -10020
rect -922 -10054 -764 -10020
rect -730 -10054 -572 -10020
rect -538 -10054 -380 -10020
rect -346 -10054 -188 -10020
rect -154 -10054 4 -10020
rect 38 -10054 196 -10020
rect 230 -10054 388 -10020
rect 422 -10054 580 -10020
rect 614 -10054 772 -10020
rect 806 -10054 964 -10020
rect 998 -10054 1156 -10020
rect 1190 -10054 1380 -10020
rect -1346 -10057 1380 -10054
rect -1346 -10060 -1102 -10057
rect -968 -10060 -910 -10057
rect -776 -10060 -718 -10057
rect -584 -10060 -526 -10057
rect -392 -10060 -334 -10057
rect -200 -10060 -142 -10057
rect -8 -10060 50 -10057
rect 184 -10060 242 -10057
rect 376 -10060 434 -10057
rect 568 -10060 626 -10057
rect 760 -10060 818 -10057
rect 952 -10060 1010 -10057
rect 1130 -10060 1380 -10057
rect -1346 -10530 -1246 -10060
rect -1202 -10104 -1156 -10092
rect -1202 -10332 -1196 -10104
rect -1162 -10332 -1156 -10104
rect -1119 -10252 -1109 -10092
rect -1057 -10252 -1047 -10092
rect -1010 -10104 -964 -10092
rect -1215 -10492 -1205 -10332
rect -1153 -10492 -1143 -10332
rect -1106 -10480 -1100 -10252
rect -1066 -10480 -1060 -10252
rect -1010 -10332 -1004 -10104
rect -970 -10332 -964 -10104
rect -927 -10252 -917 -10092
rect -865 -10252 -855 -10092
rect -818 -10104 -772 -10092
rect -1106 -10492 -1060 -10480
rect -1023 -10492 -1013 -10332
rect -961 -10492 -951 -10332
rect -914 -10480 -908 -10252
rect -874 -10480 -868 -10252
rect -818 -10332 -812 -10104
rect -778 -10332 -772 -10104
rect -735 -10252 -725 -10092
rect -673 -10252 -663 -10092
rect -626 -10104 -580 -10092
rect -914 -10492 -868 -10480
rect -831 -10492 -821 -10332
rect -769 -10492 -759 -10332
rect -722 -10480 -716 -10252
rect -682 -10480 -676 -10252
rect -626 -10332 -620 -10104
rect -586 -10332 -580 -10104
rect -543 -10252 -533 -10092
rect -481 -10252 -471 -10092
rect -434 -10104 -388 -10092
rect -722 -10492 -676 -10480
rect -639 -10492 -629 -10332
rect -577 -10492 -567 -10332
rect -530 -10480 -524 -10252
rect -490 -10480 -484 -10252
rect -434 -10332 -428 -10104
rect -394 -10332 -388 -10104
rect -351 -10252 -341 -10092
rect -289 -10252 -279 -10092
rect -242 -10104 -196 -10092
rect -530 -10492 -484 -10480
rect -447 -10492 -437 -10332
rect -385 -10492 -375 -10332
rect -338 -10480 -332 -10252
rect -298 -10480 -292 -10252
rect -242 -10332 -236 -10104
rect -202 -10332 -196 -10104
rect -159 -10252 -149 -10092
rect -97 -10252 -87 -10092
rect -50 -10104 -4 -10092
rect -338 -10492 -292 -10480
rect -255 -10492 -245 -10332
rect -193 -10492 -183 -10332
rect -146 -10480 -140 -10252
rect -106 -10480 -100 -10252
rect -50 -10332 -44 -10104
rect -10 -10332 -4 -10104
rect 33 -10252 43 -10092
rect 95 -10252 105 -10092
rect 142 -10104 188 -10092
rect -146 -10492 -100 -10480
rect -63 -10492 -53 -10332
rect -1 -10492 9 -10332
rect 46 -10480 52 -10252
rect 86 -10480 92 -10252
rect 142 -10332 148 -10104
rect 182 -10332 188 -10104
rect 225 -10252 235 -10092
rect 287 -10252 297 -10092
rect 334 -10104 380 -10092
rect 46 -10492 92 -10480
rect 129 -10492 139 -10332
rect 191 -10492 201 -10332
rect 238 -10480 244 -10252
rect 278 -10480 284 -10252
rect 334 -10332 340 -10104
rect 374 -10332 380 -10104
rect 417 -10252 427 -10092
rect 479 -10252 489 -10092
rect 526 -10104 572 -10092
rect 238 -10492 284 -10480
rect 321 -10492 331 -10332
rect 383 -10492 393 -10332
rect 430 -10480 436 -10252
rect 470 -10480 476 -10252
rect 526 -10332 532 -10104
rect 566 -10332 572 -10104
rect 609 -10252 619 -10092
rect 671 -10252 681 -10092
rect 718 -10104 764 -10092
rect 430 -10492 476 -10480
rect 513 -10492 523 -10332
rect 575 -10492 585 -10332
rect 622 -10480 628 -10252
rect 662 -10480 668 -10252
rect 718 -10332 724 -10104
rect 758 -10332 764 -10104
rect 801 -10252 811 -10092
rect 863 -10252 873 -10092
rect 910 -10104 956 -10092
rect 622 -10492 668 -10480
rect 705 -10492 715 -10332
rect 767 -10492 777 -10332
rect 814 -10480 820 -10252
rect 854 -10480 860 -10252
rect 910 -10332 916 -10104
rect 950 -10332 956 -10104
rect 993 -10252 1003 -10092
rect 1055 -10252 1065 -10092
rect 1102 -10104 1148 -10092
rect 814 -10492 860 -10480
rect 897 -10492 907 -10332
rect 959 -10492 969 -10332
rect 1006 -10480 1012 -10252
rect 1046 -10480 1052 -10252
rect 1102 -10332 1108 -10104
rect 1142 -10332 1148 -10104
rect 1185 -10252 1195 -10092
rect 1247 -10252 1257 -10092
rect 1006 -10492 1052 -10480
rect 1089 -10492 1099 -10332
rect 1151 -10492 1161 -10332
rect 1198 -10480 1204 -10252
rect 1238 -10480 1244 -10252
rect 1198 -10492 1244 -10480
rect -1064 -10527 -1006 -10524
rect -872 -10527 -814 -10524
rect -680 -10527 -622 -10524
rect -488 -10527 -430 -10524
rect -296 -10527 -238 -10524
rect -104 -10527 -46 -10524
rect 88 -10527 146 -10524
rect 280 -10527 338 -10524
rect 472 -10527 530 -10524
rect 664 -10527 722 -10524
rect 856 -10527 914 -10524
rect 1048 -10527 1106 -10524
rect -1203 -10530 1247 -10527
rect -1346 -10564 -1052 -10530
rect -1018 -10564 -860 -10530
rect -826 -10564 -668 -10530
rect -634 -10564 -476 -10530
rect -442 -10564 -284 -10530
rect -250 -10564 -92 -10530
rect -58 -10564 100 -10530
rect 134 -10564 292 -10530
rect 326 -10564 484 -10530
rect 518 -10564 676 -10530
rect 710 -10564 868 -10530
rect 902 -10564 1060 -10530
rect 1094 -10564 1247 -10530
rect -1346 -10638 1247 -10564
rect -1346 -10672 -1052 -10638
rect -1018 -10672 -860 -10638
rect -826 -10672 -668 -10638
rect -634 -10672 -476 -10638
rect -442 -10672 -284 -10638
rect -250 -10672 -92 -10638
rect -58 -10672 100 -10638
rect 134 -10672 292 -10638
rect 326 -10672 484 -10638
rect 518 -10672 676 -10638
rect 710 -10672 868 -10638
rect 902 -10672 1060 -10638
rect 1094 -10672 1247 -10638
rect -1346 -10677 1247 -10672
rect -1346 -10680 -1186 -10677
rect -1064 -10678 -1006 -10677
rect -872 -10678 -814 -10677
rect -680 -10678 -622 -10677
rect -488 -10678 -430 -10677
rect -296 -10678 -238 -10677
rect -104 -10678 -46 -10677
rect 88 -10678 146 -10677
rect 280 -10678 338 -10677
rect 472 -10678 530 -10677
rect 664 -10678 722 -10677
rect 856 -10678 914 -10677
rect 1048 -10678 1106 -10677
rect -1346 -11150 -1246 -10680
rect -1215 -10870 -1205 -10710
rect -1153 -10870 -1143 -10710
rect -1106 -10722 -1060 -10710
rect -1202 -11098 -1196 -10870
rect -1162 -11098 -1156 -10870
rect -1106 -10950 -1100 -10722
rect -1066 -10950 -1060 -10722
rect -1023 -10870 -1013 -10710
rect -961 -10870 -951 -10710
rect -914 -10722 -868 -10710
rect -1202 -11110 -1156 -11098
rect -1119 -11110 -1109 -10950
rect -1057 -11110 -1047 -10950
rect -1010 -11098 -1004 -10870
rect -970 -11098 -964 -10870
rect -914 -10950 -908 -10722
rect -874 -10950 -868 -10722
rect -831 -10870 -821 -10710
rect -769 -10870 -759 -10710
rect -722 -10722 -676 -10710
rect -1010 -11110 -964 -11098
rect -927 -11110 -917 -10950
rect -865 -11110 -855 -10950
rect -818 -11098 -812 -10870
rect -778 -11098 -772 -10870
rect -722 -10950 -716 -10722
rect -682 -10950 -676 -10722
rect -639 -10870 -629 -10710
rect -577 -10870 -567 -10710
rect -530 -10722 -484 -10710
rect -818 -11110 -772 -11098
rect -735 -11110 -725 -10950
rect -673 -11110 -663 -10950
rect -626 -11098 -620 -10870
rect -586 -11098 -580 -10870
rect -530 -10950 -524 -10722
rect -490 -10950 -484 -10722
rect -447 -10870 -437 -10710
rect -385 -10870 -375 -10710
rect -338 -10722 -292 -10710
rect -626 -11110 -580 -11098
rect -543 -11110 -533 -10950
rect -481 -11110 -471 -10950
rect -434 -11098 -428 -10870
rect -394 -11098 -388 -10870
rect -338 -10950 -332 -10722
rect -298 -10950 -292 -10722
rect -255 -10870 -245 -10710
rect -193 -10870 -183 -10710
rect -146 -10722 -100 -10710
rect -434 -11110 -388 -11098
rect -351 -11110 -341 -10950
rect -289 -11110 -279 -10950
rect -242 -11098 -236 -10870
rect -202 -11098 -196 -10870
rect -146 -10950 -140 -10722
rect -106 -10950 -100 -10722
rect -63 -10870 -53 -10710
rect -1 -10870 9 -10710
rect 46 -10722 92 -10710
rect -242 -11110 -196 -11098
rect -159 -11110 -149 -10950
rect -97 -11110 -87 -10950
rect -50 -11098 -44 -10870
rect -10 -11098 -4 -10870
rect 46 -10950 52 -10722
rect 86 -10950 92 -10722
rect 129 -10870 139 -10710
rect 191 -10870 201 -10710
rect 238 -10722 284 -10710
rect -50 -11110 -4 -11098
rect 33 -11110 43 -10950
rect 95 -11110 105 -10950
rect 142 -11098 148 -10870
rect 182 -11098 188 -10870
rect 238 -10950 244 -10722
rect 278 -10950 284 -10722
rect 321 -10870 331 -10710
rect 383 -10870 393 -10710
rect 430 -10722 476 -10710
rect 142 -11110 188 -11098
rect 225 -11110 235 -10950
rect 287 -11110 297 -10950
rect 334 -11098 340 -10870
rect 374 -11098 380 -10870
rect 430 -10950 436 -10722
rect 470 -10950 476 -10722
rect 513 -10870 523 -10710
rect 575 -10870 585 -10710
rect 622 -10722 668 -10710
rect 334 -11110 380 -11098
rect 417 -11110 427 -10950
rect 479 -11110 489 -10950
rect 526 -11098 532 -10870
rect 566 -11098 572 -10870
rect 622 -10950 628 -10722
rect 662 -10950 668 -10722
rect 705 -10870 715 -10710
rect 767 -10870 777 -10710
rect 814 -10722 860 -10710
rect 526 -11110 572 -11098
rect 609 -11110 619 -10950
rect 671 -11110 681 -10950
rect 718 -11098 724 -10870
rect 758 -11098 764 -10870
rect 814 -10950 820 -10722
rect 854 -10950 860 -10722
rect 897 -10870 907 -10710
rect 959 -10870 969 -10710
rect 1006 -10722 1052 -10710
rect 718 -11110 764 -11098
rect 801 -11110 811 -10950
rect 863 -11110 873 -10950
rect 910 -11098 916 -10870
rect 950 -11098 956 -10870
rect 1006 -10950 1012 -10722
rect 1046 -10950 1052 -10722
rect 1089 -10870 1099 -10710
rect 1151 -10870 1161 -10710
rect 1198 -10722 1244 -10710
rect 910 -11110 956 -11098
rect 993 -11110 1003 -10950
rect 1055 -11110 1065 -10950
rect 1102 -11098 1108 -10870
rect 1142 -11098 1148 -10870
rect 1198 -10950 1204 -10722
rect 1238 -10950 1244 -10722
rect 1102 -11110 1148 -11098
rect 1185 -11110 1195 -10950
rect 1247 -11110 1257 -10950
rect 1330 -10960 1380 -10060
rect 1602 -9946 1648 -9934
rect 1602 -10898 1608 -9946
rect 1642 -10898 1648 -9946
rect 1602 -10910 1648 -10898
rect 2138 -9946 2184 -9934
rect 2138 -10898 2144 -9946
rect 2178 -10898 2184 -9946
rect 2138 -10910 2184 -10898
rect 2522 -9946 2568 -9934
rect 2522 -10898 2528 -9946
rect 2562 -10898 2568 -9946
rect 2522 -10910 2568 -10898
rect 3058 -9946 3104 -9934
rect 3058 -10898 3064 -9946
rect 3098 -10898 3104 -9946
rect 3058 -10910 3104 -10898
rect 3442 -9946 3488 -9934
rect 3442 -10898 3448 -9946
rect 3482 -10898 3488 -9946
rect 3442 -10910 3488 -10898
rect 3978 -9946 4024 -9934
rect 3978 -10898 3984 -9946
rect 4018 -10898 4024 -9946
rect 3978 -10910 4024 -10898
rect 4362 -9946 4408 -9934
rect 4362 -10898 4368 -9946
rect 4402 -10898 4408 -9946
rect 4362 -10910 4408 -10898
rect 4898 -9946 4944 -9934
rect 4898 -10898 4904 -9946
rect 4938 -10898 4944 -9946
rect 4898 -10910 4944 -10898
rect 5282 -9946 5328 -9934
rect 5282 -10898 5288 -9946
rect 5322 -10898 5328 -9946
rect 5282 -10910 5328 -10898
rect 5818 -9946 5864 -9934
rect 5818 -10898 5824 -9946
rect 5858 -10898 5864 -9946
rect 5818 -10910 5864 -10898
rect 6300 -10211 6340 -9890
rect 6380 -10070 6390 -9960
rect 6460 -10070 6470 -9960
rect 6390 -10124 6450 -10070
rect 6380 -10130 6572 -10124
rect 6380 -10164 6392 -10130
rect 6560 -10164 6572 -10130
rect 6380 -10170 6572 -10164
rect 6300 -10223 6370 -10211
rect 6300 -10299 6330 -10223
rect 6364 -10299 6370 -10223
rect 6300 -10311 6370 -10299
rect 6300 -10770 6340 -10311
rect 6420 -10352 6480 -10170
rect 6664 -10200 6766 -10188
rect 6610 -10211 6620 -10200
rect 6582 -10223 6620 -10211
rect 6582 -10299 6588 -10223
rect 6582 -10311 6620 -10299
rect 6610 -10320 6620 -10311
rect 6760 -10320 6770 -10200
rect 6664 -10332 6766 -10320
rect 6380 -10358 6572 -10352
rect 6380 -10392 6392 -10358
rect 6560 -10392 6572 -10358
rect 6380 -10398 6572 -10392
rect 6420 -10692 6480 -10398
rect 6380 -10698 6572 -10692
rect 6380 -10732 6392 -10698
rect 6560 -10732 6572 -10698
rect 6380 -10738 6572 -10732
rect 6300 -10782 6370 -10770
rect 6300 -10858 6330 -10782
rect 6364 -10858 6370 -10782
rect 6300 -10870 6370 -10858
rect 1697 -10960 2089 -10954
rect 2617 -10960 3009 -10954
rect 3537 -10960 3929 -10954
rect 4457 -10960 4849 -10954
rect 5377 -10960 5769 -10954
rect 6300 -10960 6340 -10870
rect 6420 -10902 6480 -10738
rect 6582 -10782 6628 -10770
rect 6582 -10858 6588 -10782
rect 6622 -10858 6628 -10782
rect 6582 -10870 6628 -10858
rect 6380 -10908 6572 -10902
rect 6380 -10942 6392 -10908
rect 6560 -10942 6572 -10908
rect 6380 -10948 6572 -10942
rect 1330 -10994 1709 -10960
rect 2077 -10994 2629 -10960
rect 2997 -10994 3549 -10960
rect 3917 -10994 4469 -10960
rect 4837 -10994 5389 -10960
rect 5757 -10994 6340 -10960
rect 1330 -11010 6340 -10994
rect -1160 -11147 -1102 -11142
rect -968 -11147 -910 -11142
rect -776 -11147 -718 -11142
rect -584 -11147 -526 -11142
rect -392 -11147 -334 -11142
rect -200 -11147 -142 -11142
rect -8 -11147 50 -11142
rect 184 -11147 242 -11142
rect 376 -11147 434 -11142
rect 568 -11147 626 -11142
rect 760 -11147 818 -11142
rect 952 -11147 1010 -11142
rect 1144 -11147 1202 -11142
rect -1203 -11148 1247 -11147
rect -1203 -11150 -1148 -11148
rect -1346 -11182 -1148 -11150
rect -1114 -11182 -956 -11148
rect -922 -11182 -764 -11148
rect -730 -11182 -572 -11148
rect -538 -11182 -380 -11148
rect -346 -11182 -188 -11148
rect -154 -11182 4 -11148
rect 38 -11182 196 -11148
rect 230 -11182 388 -11148
rect 422 -11182 580 -11148
rect 614 -11182 772 -11148
rect 806 -11182 964 -11148
rect 998 -11182 1156 -11148
rect 1190 -11182 1247 -11148
rect -1346 -11197 1247 -11182
rect -1346 -11200 -1196 -11197
<< via1 >>
rect -1087 2533 -1035 2545
rect -1087 2385 -1078 2533
rect -1078 2385 -1044 2533
rect -1044 2385 -1035 2533
rect -1185 2157 -1176 2305
rect -1176 2157 -1142 2305
rect -1142 2157 -1133 2305
rect -1185 2145 -1133 2157
rect -891 2533 -839 2545
rect -891 2385 -882 2533
rect -882 2385 -848 2533
rect -848 2385 -839 2533
rect -989 2157 -980 2305
rect -980 2157 -946 2305
rect -946 2157 -937 2305
rect -989 2145 -937 2157
rect -695 2533 -643 2545
rect -695 2385 -686 2533
rect -686 2385 -652 2533
rect -652 2385 -643 2533
rect -793 2157 -784 2305
rect -784 2157 -750 2305
rect -750 2157 -741 2305
rect -793 2145 -741 2157
rect -499 2533 -447 2545
rect -499 2385 -490 2533
rect -490 2385 -456 2533
rect -456 2385 -447 2533
rect -597 2157 -588 2305
rect -588 2157 -554 2305
rect -554 2157 -545 2305
rect -597 2145 -545 2157
rect -303 2533 -251 2545
rect -303 2385 -294 2533
rect -294 2385 -260 2533
rect -260 2385 -251 2533
rect -401 2157 -392 2305
rect -392 2157 -358 2305
rect -358 2157 -349 2305
rect -401 2145 -349 2157
rect -107 2533 -55 2545
rect -107 2385 -98 2533
rect -98 2385 -64 2533
rect -64 2385 -55 2533
rect -205 2157 -196 2305
rect -196 2157 -162 2305
rect -162 2157 -153 2305
rect -205 2145 -153 2157
rect 89 2533 141 2545
rect 89 2385 98 2533
rect 98 2385 132 2533
rect 132 2385 141 2533
rect -9 2157 0 2305
rect 0 2157 34 2305
rect 34 2157 43 2305
rect -9 2145 43 2157
rect 285 2533 337 2545
rect 285 2385 294 2533
rect 294 2385 328 2533
rect 328 2385 337 2533
rect 187 2157 196 2305
rect 196 2157 230 2305
rect 230 2157 239 2305
rect 187 2145 239 2157
rect 711 2533 763 2545
rect 711 2385 720 2533
rect 720 2385 754 2533
rect 754 2385 763 2533
rect 613 2157 622 2305
rect 622 2157 656 2305
rect 656 2157 665 2305
rect 613 2145 665 2157
rect 907 2533 959 2545
rect 907 2385 916 2533
rect 916 2385 950 2533
rect 950 2385 959 2533
rect 809 2157 818 2305
rect 818 2157 852 2305
rect 852 2157 861 2305
rect 809 2145 861 2157
rect 1103 2533 1155 2545
rect 1103 2385 1112 2533
rect 1112 2385 1146 2533
rect 1146 2385 1155 2533
rect 1005 2157 1014 2305
rect 1014 2157 1048 2305
rect 1048 2157 1057 2305
rect 1005 2145 1057 2157
rect 1299 2533 1351 2545
rect 1299 2385 1308 2533
rect 1308 2385 1342 2533
rect 1342 2385 1351 2533
rect 1201 2157 1210 2305
rect 1210 2157 1244 2305
rect 1244 2157 1253 2305
rect 1201 2145 1253 2157
rect 1495 2533 1547 2545
rect 1495 2385 1504 2533
rect 1504 2385 1538 2533
rect 1538 2385 1547 2533
rect 1397 2157 1406 2305
rect 1406 2157 1440 2305
rect 1440 2157 1449 2305
rect 1397 2145 1449 2157
rect 1691 2533 1743 2545
rect 1691 2385 1700 2533
rect 1700 2385 1734 2533
rect 1734 2385 1743 2533
rect 1593 2157 1602 2305
rect 1602 2157 1636 2305
rect 1636 2157 1645 2305
rect 1593 2145 1645 2157
rect 1887 2533 1939 2545
rect 1887 2385 1896 2533
rect 1896 2385 1930 2533
rect 1930 2385 1939 2533
rect 1789 2157 1798 2305
rect 1798 2157 1832 2305
rect 1832 2157 1841 2305
rect 1789 2145 1841 2157
rect 2083 2533 2135 2545
rect 2083 2385 2092 2533
rect 2092 2385 2126 2533
rect 2126 2385 2135 2533
rect 1985 2157 1994 2305
rect 1994 2157 2028 2305
rect 2028 2157 2037 2305
rect 1985 2145 2037 2157
rect -1185 1897 -1133 1909
rect -1185 1749 -1176 1897
rect -1176 1749 -1142 1897
rect -1142 1749 -1133 1897
rect -989 1897 -937 1909
rect -989 1749 -980 1897
rect -980 1749 -946 1897
rect -946 1749 -937 1897
rect -1087 1521 -1078 1669
rect -1078 1521 -1044 1669
rect -1044 1521 -1035 1669
rect -1087 1509 -1035 1521
rect -793 1897 -741 1909
rect -793 1749 -784 1897
rect -784 1749 -750 1897
rect -750 1749 -741 1897
rect -891 1521 -882 1669
rect -882 1521 -848 1669
rect -848 1521 -839 1669
rect -891 1509 -839 1521
rect -597 1897 -545 1909
rect -597 1749 -588 1897
rect -588 1749 -554 1897
rect -554 1749 -545 1897
rect -695 1521 -686 1669
rect -686 1521 -652 1669
rect -652 1521 -643 1669
rect -695 1509 -643 1521
rect -401 1897 -349 1909
rect -401 1749 -392 1897
rect -392 1749 -358 1897
rect -358 1749 -349 1897
rect -499 1521 -490 1669
rect -490 1521 -456 1669
rect -456 1521 -447 1669
rect -499 1509 -447 1521
rect -205 1897 -153 1909
rect -205 1749 -196 1897
rect -196 1749 -162 1897
rect -162 1749 -153 1897
rect -303 1521 -294 1669
rect -294 1521 -260 1669
rect -260 1521 -251 1669
rect -303 1509 -251 1521
rect -9 1897 43 1909
rect -9 1749 0 1897
rect 0 1749 34 1897
rect 34 1749 43 1897
rect -107 1521 -98 1669
rect -98 1521 -64 1669
rect -64 1521 -55 1669
rect -107 1509 -55 1521
rect 187 1897 239 1909
rect 187 1749 196 1897
rect 196 1749 230 1897
rect 230 1749 239 1897
rect 89 1521 98 1669
rect 98 1521 132 1669
rect 132 1521 141 1669
rect 89 1509 141 1521
rect 285 1521 294 1669
rect 294 1521 328 1669
rect 328 1521 337 1669
rect 285 1509 337 1521
rect 613 1897 665 1909
rect 613 1749 622 1897
rect 622 1749 656 1897
rect 656 1749 665 1897
rect 809 1897 861 1909
rect 809 1749 818 1897
rect 818 1749 852 1897
rect 852 1749 861 1897
rect 711 1521 720 1669
rect 720 1521 754 1669
rect 754 1521 763 1669
rect 711 1509 763 1521
rect 1005 1897 1057 1909
rect 1005 1749 1014 1897
rect 1014 1749 1048 1897
rect 1048 1749 1057 1897
rect 907 1521 916 1669
rect 916 1521 950 1669
rect 950 1521 959 1669
rect 907 1509 959 1521
rect 1201 1897 1253 1909
rect 1201 1749 1210 1897
rect 1210 1749 1244 1897
rect 1244 1749 1253 1897
rect 1103 1521 1112 1669
rect 1112 1521 1146 1669
rect 1146 1521 1155 1669
rect 1103 1509 1155 1521
rect 1397 1897 1449 1909
rect 1397 1749 1406 1897
rect 1406 1749 1440 1897
rect 1440 1749 1449 1897
rect 1299 1521 1308 1669
rect 1308 1521 1342 1669
rect 1342 1521 1351 1669
rect 1299 1509 1351 1521
rect 1593 1897 1645 1909
rect 1593 1749 1602 1897
rect 1602 1749 1636 1897
rect 1636 1749 1645 1897
rect 1495 1521 1504 1669
rect 1504 1521 1538 1669
rect 1538 1521 1547 1669
rect 1495 1509 1547 1521
rect 1789 1897 1841 1909
rect 1789 1749 1798 1897
rect 1798 1749 1832 1897
rect 1832 1749 1841 1897
rect 1691 1521 1700 1669
rect 1700 1521 1734 1669
rect 1734 1521 1743 1669
rect 1691 1509 1743 1521
rect 1985 1897 2037 1909
rect 1985 1749 1994 1897
rect 1994 1749 2028 1897
rect 2028 1749 2037 1897
rect 1887 1521 1896 1669
rect 1896 1521 1930 1669
rect 1930 1521 1939 1669
rect 1887 1509 1939 1521
rect 2083 1521 2092 1669
rect 2092 1521 2126 1669
rect 2126 1521 2135 1669
rect 2083 1509 2135 1521
rect 2214 1510 2344 2070
rect 4660 1930 4740 2000
rect 2573 1881 2625 1893
rect 2573 1733 2582 1881
rect 2582 1733 2616 1881
rect 2616 1733 2625 1881
rect 2415 1505 2424 1653
rect 2424 1505 2458 1653
rect 2458 1505 2467 1653
rect 2415 1493 2467 1505
rect 2889 1881 2941 1893
rect 2889 1733 2898 1881
rect 2898 1733 2932 1881
rect 2932 1733 2941 1881
rect 2731 1505 2740 1653
rect 2740 1505 2774 1653
rect 2774 1505 2783 1653
rect 2731 1493 2783 1505
rect 3205 1881 3257 1893
rect 3205 1733 3214 1881
rect 3214 1733 3248 1881
rect 3248 1733 3257 1881
rect 3047 1505 3056 1653
rect 3056 1505 3090 1653
rect 3090 1505 3099 1653
rect 3047 1493 3099 1505
rect 3521 1881 3573 1893
rect 3521 1733 3530 1881
rect 3530 1733 3564 1881
rect 3564 1733 3573 1881
rect 3363 1505 3372 1653
rect 3372 1505 3406 1653
rect 3406 1505 3415 1653
rect 3363 1493 3415 1505
rect 3837 1881 3889 1893
rect 3837 1733 3846 1881
rect 3846 1733 3880 1881
rect 3880 1733 3889 1881
rect 3679 1505 3688 1653
rect 3688 1505 3722 1653
rect 3722 1505 3731 1653
rect 3679 1493 3731 1505
rect 3995 1505 4004 1653
rect 4004 1505 4038 1653
rect 4038 1505 4047 1653
rect 3995 1493 4047 1505
rect -1087 1066 -1035 1078
rect -1087 918 -1078 1066
rect -1078 918 -1044 1066
rect -1044 918 -1035 1066
rect -1185 690 -1176 838
rect -1176 690 -1142 838
rect -1142 690 -1133 838
rect -1185 678 -1133 690
rect -891 1066 -839 1078
rect -891 918 -882 1066
rect -882 918 -848 1066
rect -848 918 -839 1066
rect -989 690 -980 838
rect -980 690 -946 838
rect -946 690 -937 838
rect -989 678 -937 690
rect -695 1066 -643 1078
rect -695 918 -686 1066
rect -686 918 -652 1066
rect -652 918 -643 1066
rect -793 690 -784 838
rect -784 690 -750 838
rect -750 690 -741 838
rect -793 678 -741 690
rect -499 1066 -447 1078
rect -499 918 -490 1066
rect -490 918 -456 1066
rect -456 918 -447 1066
rect -597 690 -588 838
rect -588 690 -554 838
rect -554 690 -545 838
rect -597 678 -545 690
rect -303 1066 -251 1078
rect -303 918 -294 1066
rect -294 918 -260 1066
rect -260 918 -251 1066
rect -401 690 -392 838
rect -392 690 -358 838
rect -358 690 -349 838
rect -401 678 -349 690
rect -107 1066 -55 1078
rect -107 918 -98 1066
rect -98 918 -64 1066
rect -64 918 -55 1066
rect -205 690 -196 838
rect -196 690 -162 838
rect -162 690 -153 838
rect -205 678 -153 690
rect 89 1066 141 1078
rect 89 918 98 1066
rect 98 918 132 1066
rect 132 918 141 1066
rect -9 690 0 838
rect 0 690 34 838
rect 34 690 43 838
rect -9 678 43 690
rect 285 1066 337 1078
rect 285 918 294 1066
rect 294 918 328 1066
rect 328 918 337 1066
rect 187 690 196 838
rect 196 690 230 838
rect 230 690 239 838
rect 187 678 239 690
rect 481 1066 533 1078
rect 481 918 490 1066
rect 490 918 524 1066
rect 524 918 533 1066
rect 383 690 392 838
rect 392 690 426 838
rect 426 690 435 838
rect 383 678 435 690
rect 677 1066 729 1078
rect 677 918 686 1066
rect 686 918 720 1066
rect 720 918 729 1066
rect 579 690 588 838
rect 588 690 622 838
rect 622 690 631 838
rect 579 678 631 690
rect 873 1066 925 1078
rect 873 918 882 1066
rect 882 918 916 1066
rect 916 918 925 1066
rect 775 690 784 838
rect 784 690 818 838
rect 818 690 827 838
rect 775 678 827 690
rect 1069 1066 1121 1078
rect 1069 918 1078 1066
rect 1078 918 1112 1066
rect 1112 918 1121 1066
rect 971 690 980 838
rect 980 690 1014 838
rect 1014 690 1023 838
rect 971 678 1023 690
rect 1265 1066 1317 1078
rect 1265 918 1274 1066
rect 1274 918 1308 1066
rect 1308 918 1317 1066
rect 1167 690 1176 838
rect 1176 690 1210 838
rect 1210 690 1219 838
rect 1167 678 1219 690
rect 2164 660 2414 850
rect -1185 448 -1133 460
rect -1185 300 -1176 448
rect -1176 300 -1142 448
rect -1142 300 -1133 448
rect -989 448 -937 460
rect -989 300 -980 448
rect -980 300 -946 448
rect -946 300 -937 448
rect -1087 72 -1078 220
rect -1078 72 -1044 220
rect -1044 72 -1035 220
rect -1087 60 -1035 72
rect -793 448 -741 460
rect -793 300 -784 448
rect -784 300 -750 448
rect -750 300 -741 448
rect -891 72 -882 220
rect -882 72 -848 220
rect -848 72 -839 220
rect -891 60 -839 72
rect -597 448 -545 460
rect -597 300 -588 448
rect -588 300 -554 448
rect -554 300 -545 448
rect -695 72 -686 220
rect -686 72 -652 220
rect -652 72 -643 220
rect -695 60 -643 72
rect -401 448 -349 460
rect -401 300 -392 448
rect -392 300 -358 448
rect -358 300 -349 448
rect -499 72 -490 220
rect -490 72 -456 220
rect -456 72 -447 220
rect -499 60 -447 72
rect -205 448 -153 460
rect -205 300 -196 448
rect -196 300 -162 448
rect -162 300 -153 448
rect -303 72 -294 220
rect -294 72 -260 220
rect -260 72 -251 220
rect -303 60 -251 72
rect -9 448 43 460
rect -9 300 0 448
rect 0 300 34 448
rect 34 300 43 448
rect -107 72 -98 220
rect -98 72 -64 220
rect -64 72 -55 220
rect -107 60 -55 72
rect 187 448 239 460
rect 187 300 196 448
rect 196 300 230 448
rect 230 300 239 448
rect 89 72 98 220
rect 98 72 132 220
rect 132 72 141 220
rect 89 60 141 72
rect 383 448 435 460
rect 383 300 392 448
rect 392 300 426 448
rect 426 300 435 448
rect 285 72 294 220
rect 294 72 328 220
rect 328 72 337 220
rect 285 60 337 72
rect 579 448 631 460
rect 579 300 588 448
rect 588 300 622 448
rect 622 300 631 448
rect 481 72 490 220
rect 490 72 524 220
rect 524 72 533 220
rect 481 60 533 72
rect 775 448 827 460
rect 775 300 784 448
rect 784 300 818 448
rect 818 300 827 448
rect 677 72 686 220
rect 686 72 720 220
rect 720 72 729 220
rect 677 60 729 72
rect 971 448 1023 460
rect 971 300 980 448
rect 980 300 1014 448
rect 1014 300 1023 448
rect 873 72 882 220
rect 882 72 916 220
rect 916 72 925 220
rect 873 60 925 72
rect 1167 448 1219 460
rect 1167 300 1176 448
rect 1176 300 1210 448
rect 1210 300 1219 448
rect 1069 72 1078 220
rect 1078 72 1112 220
rect 1112 72 1121 220
rect 1069 60 1121 72
rect 2475 746 2527 758
rect 2475 598 2484 746
rect 2484 598 2518 746
rect 2518 598 2527 746
rect 2671 746 2723 758
rect 2671 598 2680 746
rect 2680 598 2714 746
rect 2714 598 2723 746
rect 2573 370 2582 518
rect 2582 370 2616 518
rect 2616 370 2625 518
rect 2573 358 2625 370
rect 2867 746 2919 758
rect 2867 598 2876 746
rect 2876 598 2910 746
rect 2910 598 2919 746
rect 2769 370 2778 518
rect 2778 370 2812 518
rect 2812 370 2821 518
rect 2769 358 2821 370
rect 3063 746 3115 758
rect 3063 598 3072 746
rect 3072 598 3106 746
rect 3106 598 3115 746
rect 2965 370 2974 518
rect 2974 370 3008 518
rect 3008 370 3017 518
rect 2965 358 3017 370
rect 3259 746 3311 758
rect 3259 598 3268 746
rect 3268 598 3302 746
rect 3302 598 3311 746
rect 3161 370 3170 518
rect 3170 370 3204 518
rect 3204 370 3213 518
rect 3161 358 3213 370
rect 3455 746 3507 758
rect 3455 598 3464 746
rect 3464 598 3498 746
rect 3498 598 3507 746
rect 3357 370 3366 518
rect 3366 370 3400 518
rect 3400 370 3409 518
rect 3357 358 3409 370
rect 3651 746 3703 758
rect 3651 598 3660 746
rect 3660 598 3694 746
rect 3694 598 3703 746
rect 3553 370 3562 518
rect 3562 370 3596 518
rect 3596 370 3605 518
rect 3553 358 3605 370
rect 3847 746 3899 758
rect 3847 598 3856 746
rect 3856 598 3890 746
rect 3890 598 3899 746
rect 3749 370 3758 518
rect 3758 370 3792 518
rect 3792 370 3801 518
rect 3749 358 3801 370
rect 3945 370 3954 518
rect 3954 370 3988 518
rect 3988 370 3997 518
rect 3945 358 3997 370
rect 1265 72 1274 220
rect 1274 72 1308 220
rect 1308 72 1317 220
rect 1265 60 1317 72
rect 1454 160 1684 320
rect 2204 160 2284 320
rect -1087 -378 -1035 -366
rect -1087 -526 -1078 -378
rect -1078 -526 -1044 -378
rect -1044 -526 -1035 -378
rect -1185 -754 -1176 -606
rect -1176 -754 -1142 -606
rect -1142 -754 -1133 -606
rect -1185 -766 -1133 -754
rect -891 -378 -839 -366
rect -891 -526 -882 -378
rect -882 -526 -848 -378
rect -848 -526 -839 -378
rect -989 -754 -980 -606
rect -980 -754 -946 -606
rect -946 -754 -937 -606
rect -989 -766 -937 -754
rect -695 -378 -643 -366
rect -695 -526 -686 -378
rect -686 -526 -652 -378
rect -652 -526 -643 -378
rect -793 -754 -784 -606
rect -784 -754 -750 -606
rect -750 -754 -741 -606
rect -793 -766 -741 -754
rect -499 -378 -447 -366
rect -499 -526 -490 -378
rect -490 -526 -456 -378
rect -456 -526 -447 -378
rect -597 -754 -588 -606
rect -588 -754 -554 -606
rect -554 -754 -545 -606
rect -597 -766 -545 -754
rect -303 -378 -251 -366
rect -303 -526 -294 -378
rect -294 -526 -260 -378
rect -260 -526 -251 -378
rect -401 -754 -392 -606
rect -392 -754 -358 -606
rect -358 -754 -349 -606
rect -401 -766 -349 -754
rect -107 -378 -55 -366
rect -107 -526 -98 -378
rect -98 -526 -64 -378
rect -64 -526 -55 -378
rect -205 -754 -196 -606
rect -196 -754 -162 -606
rect -162 -754 -153 -606
rect -205 -766 -153 -754
rect 89 -378 141 -366
rect 89 -526 98 -378
rect 98 -526 132 -378
rect 132 -526 141 -378
rect -9 -754 0 -606
rect 0 -754 34 -606
rect 34 -754 43 -606
rect -9 -766 43 -754
rect 285 -378 337 -366
rect 285 -526 294 -378
rect 294 -526 328 -378
rect 328 -526 337 -378
rect 187 -754 196 -606
rect 196 -754 230 -606
rect 230 -754 239 -606
rect 187 -766 239 -754
rect 481 -378 533 -366
rect 481 -526 490 -378
rect 490 -526 524 -378
rect 524 -526 533 -378
rect 383 -754 392 -606
rect 392 -754 426 -606
rect 426 -754 435 -606
rect 383 -766 435 -754
rect 677 -378 729 -366
rect 677 -526 686 -378
rect 686 -526 720 -378
rect 720 -526 729 -378
rect 579 -754 588 -606
rect 588 -754 622 -606
rect 622 -754 631 -606
rect 579 -766 631 -754
rect 873 -378 925 -366
rect 873 -526 882 -378
rect 882 -526 916 -378
rect 916 -526 925 -378
rect 775 -754 784 -606
rect 784 -754 818 -606
rect 818 -754 827 -606
rect 775 -766 827 -754
rect 1069 -378 1121 -366
rect 1069 -526 1078 -378
rect 1078 -526 1112 -378
rect 1112 -526 1121 -378
rect 971 -754 980 -606
rect 980 -754 1014 -606
rect 1014 -754 1023 -606
rect 971 -766 1023 -754
rect 1265 -378 1317 -366
rect 1265 -526 1274 -378
rect 1274 -526 1308 -378
rect 1308 -526 1317 -378
rect 1167 -754 1176 -606
rect 1176 -754 1210 -606
rect 1210 -754 1219 -606
rect 1167 -766 1219 -754
rect 2573 128 2625 140
rect 2573 -20 2582 128
rect 2582 -20 2616 128
rect 2616 -20 2625 128
rect 2475 -248 2484 -100
rect 2484 -248 2518 -100
rect 2518 -248 2527 -100
rect 2475 -260 2527 -248
rect 2769 128 2821 140
rect 2769 -20 2778 128
rect 2778 -20 2812 128
rect 2812 -20 2821 128
rect 2671 -248 2680 -100
rect 2680 -248 2714 -100
rect 2714 -248 2723 -100
rect 2671 -260 2723 -248
rect 2965 128 3017 140
rect 2965 -20 2974 128
rect 2974 -20 3008 128
rect 3008 -20 3017 128
rect 2867 -248 2876 -100
rect 2876 -248 2910 -100
rect 2910 -248 2919 -100
rect 2867 -260 2919 -248
rect 3161 128 3213 140
rect 3161 -20 3170 128
rect 3170 -20 3204 128
rect 3204 -20 3213 128
rect 3063 -248 3072 -100
rect 3072 -248 3106 -100
rect 3106 -248 3115 -100
rect 3063 -260 3115 -248
rect 3357 128 3409 140
rect 3357 -20 3366 128
rect 3366 -20 3400 128
rect 3400 -20 3409 128
rect 3259 -248 3268 -100
rect 3268 -248 3302 -100
rect 3302 -248 3311 -100
rect 3259 -260 3311 -248
rect 3553 128 3605 140
rect 3553 -20 3562 128
rect 3562 -20 3596 128
rect 3596 -20 3605 128
rect 3455 -248 3464 -100
rect 3464 -248 3498 -100
rect 3498 -248 3507 -100
rect 3455 -260 3507 -248
rect 3749 128 3801 140
rect 3749 -20 3758 128
rect 3758 -20 3792 128
rect 3792 -20 3801 128
rect 3651 -248 3660 -100
rect 3660 -248 3694 -100
rect 3694 -248 3703 -100
rect 3651 -260 3703 -248
rect 3945 128 3997 140
rect 3945 -20 3954 128
rect 3954 -20 3988 128
rect 3988 -20 3997 128
rect 4054 130 4174 340
rect 3847 -248 3856 -100
rect 3856 -248 3890 -100
rect 3890 -248 3899 -100
rect 3847 -260 3899 -248
rect -1185 -996 -1133 -984
rect -1185 -1144 -1176 -996
rect -1176 -1144 -1142 -996
rect -1142 -1144 -1133 -996
rect -989 -996 -937 -984
rect -989 -1144 -980 -996
rect -980 -1144 -946 -996
rect -946 -1144 -937 -996
rect -1087 -1372 -1078 -1224
rect -1078 -1372 -1044 -1224
rect -1044 -1372 -1035 -1224
rect -1087 -1384 -1035 -1372
rect -793 -996 -741 -984
rect -793 -1144 -784 -996
rect -784 -1144 -750 -996
rect -750 -1144 -741 -996
rect -891 -1372 -882 -1224
rect -882 -1372 -848 -1224
rect -848 -1372 -839 -1224
rect -891 -1384 -839 -1372
rect -597 -996 -545 -984
rect -597 -1144 -588 -996
rect -588 -1144 -554 -996
rect -554 -1144 -545 -996
rect -695 -1372 -686 -1224
rect -686 -1372 -652 -1224
rect -652 -1372 -643 -1224
rect -695 -1384 -643 -1372
rect -401 -996 -349 -984
rect -401 -1144 -392 -996
rect -392 -1144 -358 -996
rect -358 -1144 -349 -996
rect -499 -1372 -490 -1224
rect -490 -1372 -456 -1224
rect -456 -1372 -447 -1224
rect -499 -1384 -447 -1372
rect -205 -996 -153 -984
rect -205 -1144 -196 -996
rect -196 -1144 -162 -996
rect -162 -1144 -153 -996
rect -303 -1372 -294 -1224
rect -294 -1372 -260 -1224
rect -260 -1372 -251 -1224
rect -303 -1384 -251 -1372
rect -9 -996 43 -984
rect -9 -1144 0 -996
rect 0 -1144 34 -996
rect 34 -1144 43 -996
rect -107 -1372 -98 -1224
rect -98 -1372 -64 -1224
rect -64 -1372 -55 -1224
rect -107 -1384 -55 -1372
rect 187 -996 239 -984
rect 187 -1144 196 -996
rect 196 -1144 230 -996
rect 230 -1144 239 -996
rect 89 -1372 98 -1224
rect 98 -1372 132 -1224
rect 132 -1372 141 -1224
rect 89 -1384 141 -1372
rect 383 -996 435 -984
rect 383 -1144 392 -996
rect 392 -1144 426 -996
rect 426 -1144 435 -996
rect 285 -1372 294 -1224
rect 294 -1372 328 -1224
rect 328 -1372 337 -1224
rect 285 -1384 337 -1372
rect 579 -996 631 -984
rect 579 -1144 588 -996
rect 588 -1144 622 -996
rect 622 -1144 631 -996
rect 481 -1372 490 -1224
rect 490 -1372 524 -1224
rect 524 -1372 533 -1224
rect 481 -1384 533 -1372
rect 775 -996 827 -984
rect 775 -1144 784 -996
rect 784 -1144 818 -996
rect 818 -1144 827 -996
rect 677 -1372 686 -1224
rect 686 -1372 720 -1224
rect 720 -1372 729 -1224
rect 677 -1384 729 -1372
rect 971 -996 1023 -984
rect 971 -1144 980 -996
rect 980 -1144 1014 -996
rect 1014 -1144 1023 -996
rect 873 -1372 882 -1224
rect 882 -1372 916 -1224
rect 916 -1372 925 -1224
rect 873 -1384 925 -1372
rect 1167 -996 1219 -984
rect 1167 -1144 1176 -996
rect 1176 -1144 1210 -996
rect 1210 -1144 1219 -996
rect 1069 -1372 1078 -1224
rect 1078 -1372 1112 -1224
rect 1112 -1372 1121 -1224
rect 1069 -1384 1121 -1372
rect 1265 -1372 1274 -1224
rect 1274 -1372 1308 -1224
rect 1308 -1372 1317 -1224
rect 1265 -1384 1317 -1372
rect 1701 -1032 1753 -1020
rect 1701 -1180 1710 -1032
rect 1710 -1180 1744 -1032
rect 1744 -1180 1753 -1032
rect 1605 -1408 1614 -1260
rect 1614 -1408 1648 -1260
rect 1648 -1408 1657 -1260
rect 1605 -1420 1657 -1408
rect 1893 -1032 1945 -1020
rect 1893 -1180 1902 -1032
rect 1902 -1180 1936 -1032
rect 1936 -1180 1945 -1032
rect 1797 -1408 1806 -1260
rect 1806 -1408 1840 -1260
rect 1840 -1408 1849 -1260
rect 1797 -1420 1849 -1408
rect 2085 -1032 2137 -1020
rect 2085 -1180 2094 -1032
rect 2094 -1180 2128 -1032
rect 2128 -1180 2137 -1032
rect 1989 -1408 1998 -1260
rect 1998 -1408 2032 -1260
rect 2032 -1408 2041 -1260
rect 1989 -1420 2041 -1408
rect 2277 -1032 2329 -1020
rect 2277 -1180 2286 -1032
rect 2286 -1180 2320 -1032
rect 2320 -1180 2329 -1032
rect 2181 -1408 2190 -1260
rect 2190 -1408 2224 -1260
rect 2224 -1408 2233 -1260
rect 2181 -1420 2233 -1408
rect 2469 -1032 2521 -1020
rect 2469 -1180 2478 -1032
rect 2478 -1180 2512 -1032
rect 2512 -1180 2521 -1032
rect 2373 -1408 2382 -1260
rect 2382 -1408 2416 -1260
rect 2416 -1408 2425 -1260
rect 2373 -1420 2425 -1408
rect 2661 -1032 2713 -1020
rect 2661 -1180 2670 -1032
rect 2670 -1180 2704 -1032
rect 2704 -1180 2713 -1032
rect 2565 -1408 2574 -1260
rect 2574 -1408 2608 -1260
rect 2608 -1408 2617 -1260
rect 2565 -1420 2617 -1408
rect 2757 -1408 2766 -1260
rect 2766 -1408 2800 -1260
rect 2800 -1408 2809 -1260
rect 2757 -1420 2809 -1408
rect -1109 -1798 -1057 -1786
rect -1109 -1946 -1100 -1798
rect -1100 -1946 -1066 -1798
rect -1066 -1946 -1057 -1798
rect -1205 -2174 -1196 -2026
rect -1196 -2174 -1162 -2026
rect -1162 -2174 -1153 -2026
rect -1205 -2186 -1153 -2174
rect -917 -1798 -865 -1786
rect -917 -1946 -908 -1798
rect -908 -1946 -874 -1798
rect -874 -1946 -865 -1798
rect -1013 -2174 -1004 -2026
rect -1004 -2174 -970 -2026
rect -970 -2174 -961 -2026
rect -1013 -2186 -961 -2174
rect -725 -1798 -673 -1786
rect -725 -1946 -716 -1798
rect -716 -1946 -682 -1798
rect -682 -1946 -673 -1798
rect -821 -2174 -812 -2026
rect -812 -2174 -778 -2026
rect -778 -2174 -769 -2026
rect -821 -2186 -769 -2174
rect -533 -1798 -481 -1786
rect -533 -1946 -524 -1798
rect -524 -1946 -490 -1798
rect -490 -1946 -481 -1798
rect -629 -2174 -620 -2026
rect -620 -2174 -586 -2026
rect -586 -2174 -577 -2026
rect -629 -2186 -577 -2174
rect -341 -1798 -289 -1786
rect -341 -1946 -332 -1798
rect -332 -1946 -298 -1798
rect -298 -1946 -289 -1798
rect -437 -2174 -428 -2026
rect -428 -2174 -394 -2026
rect -394 -2174 -385 -2026
rect -437 -2186 -385 -2174
rect -149 -1798 -97 -1786
rect -149 -1946 -140 -1798
rect -140 -1946 -106 -1798
rect -106 -1946 -97 -1798
rect -245 -2174 -236 -2026
rect -236 -2174 -202 -2026
rect -202 -2174 -193 -2026
rect -245 -2186 -193 -2174
rect 43 -1798 95 -1786
rect 43 -1946 52 -1798
rect 52 -1946 86 -1798
rect 86 -1946 95 -1798
rect -53 -2174 -44 -2026
rect -44 -2174 -10 -2026
rect -10 -2174 -1 -2026
rect -53 -2186 -1 -2174
rect 235 -1798 287 -1786
rect 235 -1946 244 -1798
rect 244 -1946 278 -1798
rect 278 -1946 287 -1798
rect 139 -2174 148 -2026
rect 148 -2174 182 -2026
rect 182 -2174 191 -2026
rect 139 -2186 191 -2174
rect 427 -1798 479 -1786
rect 427 -1946 436 -1798
rect 436 -1946 470 -1798
rect 470 -1946 479 -1798
rect 331 -2174 340 -2026
rect 340 -2174 374 -2026
rect 374 -2174 383 -2026
rect 331 -2186 383 -2174
rect 619 -1798 671 -1786
rect 619 -1946 628 -1798
rect 628 -1946 662 -1798
rect 662 -1946 671 -1798
rect 523 -2174 532 -2026
rect 532 -2174 566 -2026
rect 566 -2174 575 -2026
rect 523 -2186 575 -2174
rect 811 -1798 863 -1786
rect 811 -1946 820 -1798
rect 820 -1946 854 -1798
rect 854 -1946 863 -1798
rect 715 -2174 724 -2026
rect 724 -2174 758 -2026
rect 758 -2174 767 -2026
rect 715 -2186 767 -2174
rect 1003 -1798 1055 -1786
rect 1003 -1946 1012 -1798
rect 1012 -1946 1046 -1798
rect 1046 -1946 1055 -1798
rect 907 -2174 916 -2026
rect 916 -2174 950 -2026
rect 950 -2174 959 -2026
rect 907 -2186 959 -2174
rect 1195 -1798 1247 -1786
rect 1195 -1946 1204 -1798
rect 1204 -1946 1238 -1798
rect 1238 -1946 1247 -1798
rect 3140 -1780 3320 -1660
rect 1099 -2174 1108 -2026
rect 1108 -2174 1142 -2026
rect 1142 -2174 1151 -2026
rect 1099 -2186 1151 -2174
rect 1344 -2250 1474 -2070
rect 1863 -1852 1915 -1840
rect 1863 -2000 1872 -1852
rect 1872 -2000 1906 -1852
rect 1906 -2000 1915 -1852
rect 1605 -2228 1614 -2080
rect 1614 -2228 1648 -2080
rect 1648 -2228 1657 -2080
rect 1605 -2240 1657 -2228
rect 2379 -1852 2431 -1840
rect 2379 -2000 2388 -1852
rect 2388 -2000 2422 -1852
rect 2422 -2000 2431 -1852
rect 2121 -2228 2130 -2080
rect 2130 -2228 2164 -2080
rect 2164 -2228 2173 -2080
rect 2121 -2240 2173 -2228
rect 2895 -1852 2947 -1840
rect 2895 -2000 2904 -1852
rect 2904 -2000 2938 -1852
rect 2938 -2000 2947 -1852
rect 2637 -2228 2646 -2080
rect 2646 -2228 2680 -2080
rect 2680 -2228 2689 -2080
rect 2637 -2240 2689 -2228
rect 3153 -2228 3162 -2080
rect 3162 -2228 3196 -2080
rect 3196 -2228 3205 -2080
rect 3153 -2240 3205 -2228
rect -1205 -2416 -1153 -2404
rect -1205 -2564 -1196 -2416
rect -1196 -2564 -1162 -2416
rect -1162 -2564 -1153 -2416
rect -1013 -2416 -961 -2404
rect -1013 -2564 -1004 -2416
rect -1004 -2564 -970 -2416
rect -970 -2564 -961 -2416
rect -1109 -2792 -1100 -2644
rect -1100 -2792 -1066 -2644
rect -1066 -2792 -1057 -2644
rect -1109 -2804 -1057 -2792
rect -821 -2416 -769 -2404
rect -821 -2564 -812 -2416
rect -812 -2564 -778 -2416
rect -778 -2564 -769 -2416
rect -917 -2792 -908 -2644
rect -908 -2792 -874 -2644
rect -874 -2792 -865 -2644
rect -917 -2804 -865 -2792
rect -629 -2416 -577 -2404
rect -629 -2564 -620 -2416
rect -620 -2564 -586 -2416
rect -586 -2564 -577 -2416
rect -725 -2792 -716 -2644
rect -716 -2792 -682 -2644
rect -682 -2792 -673 -2644
rect -725 -2804 -673 -2792
rect -437 -2416 -385 -2404
rect -437 -2564 -428 -2416
rect -428 -2564 -394 -2416
rect -394 -2564 -385 -2416
rect -533 -2792 -524 -2644
rect -524 -2792 -490 -2644
rect -490 -2792 -481 -2644
rect -533 -2804 -481 -2792
rect -245 -2416 -193 -2404
rect -245 -2564 -236 -2416
rect -236 -2564 -202 -2416
rect -202 -2564 -193 -2416
rect -341 -2792 -332 -2644
rect -332 -2792 -298 -2644
rect -298 -2792 -289 -2644
rect -341 -2804 -289 -2792
rect -53 -2416 -1 -2404
rect -53 -2564 -44 -2416
rect -44 -2564 -10 -2416
rect -10 -2564 -1 -2416
rect -149 -2792 -140 -2644
rect -140 -2792 -106 -2644
rect -106 -2792 -97 -2644
rect -149 -2804 -97 -2792
rect 139 -2416 191 -2404
rect 139 -2564 148 -2416
rect 148 -2564 182 -2416
rect 182 -2564 191 -2416
rect 43 -2792 52 -2644
rect 52 -2792 86 -2644
rect 86 -2792 95 -2644
rect 43 -2804 95 -2792
rect 331 -2416 383 -2404
rect 331 -2564 340 -2416
rect 340 -2564 374 -2416
rect 374 -2564 383 -2416
rect 235 -2792 244 -2644
rect 244 -2792 278 -2644
rect 278 -2792 287 -2644
rect 235 -2804 287 -2792
rect 523 -2416 575 -2404
rect 523 -2564 532 -2416
rect 532 -2564 566 -2416
rect 566 -2564 575 -2416
rect 427 -2792 436 -2644
rect 436 -2792 470 -2644
rect 470 -2792 479 -2644
rect 427 -2804 479 -2792
rect 715 -2416 767 -2404
rect 715 -2564 724 -2416
rect 724 -2564 758 -2416
rect 758 -2564 767 -2416
rect 619 -2792 628 -2644
rect 628 -2792 662 -2644
rect 662 -2792 671 -2644
rect 619 -2804 671 -2792
rect 907 -2416 959 -2404
rect 907 -2564 916 -2416
rect 916 -2564 950 -2416
rect 950 -2564 959 -2416
rect 811 -2792 820 -2644
rect 820 -2792 854 -2644
rect 854 -2792 863 -2644
rect 811 -2804 863 -2792
rect 1099 -2416 1151 -2404
rect 1099 -2564 1108 -2416
rect 1108 -2564 1142 -2416
rect 1142 -2564 1151 -2416
rect 1003 -2792 1012 -2644
rect 1012 -2792 1046 -2644
rect 1046 -2792 1055 -2644
rect 1003 -2804 1055 -2792
rect 1195 -2792 1204 -2644
rect 1204 -2792 1238 -2644
rect 1238 -2792 1247 -2644
rect 1195 -2804 1247 -2792
rect -1109 -3034 -1057 -3022
rect -1109 -3182 -1100 -3034
rect -1100 -3182 -1066 -3034
rect -1066 -3182 -1057 -3034
rect -1205 -3410 -1196 -3262
rect -1196 -3410 -1162 -3262
rect -1162 -3410 -1153 -3262
rect -1205 -3422 -1153 -3410
rect -917 -3034 -865 -3022
rect -917 -3182 -908 -3034
rect -908 -3182 -874 -3034
rect -874 -3182 -865 -3034
rect -1013 -3410 -1004 -3262
rect -1004 -3410 -970 -3262
rect -970 -3410 -961 -3262
rect -1013 -3422 -961 -3410
rect -725 -3034 -673 -3022
rect -725 -3182 -716 -3034
rect -716 -3182 -682 -3034
rect -682 -3182 -673 -3034
rect -821 -3410 -812 -3262
rect -812 -3410 -778 -3262
rect -778 -3410 -769 -3262
rect -821 -3422 -769 -3410
rect -533 -3034 -481 -3022
rect -533 -3182 -524 -3034
rect -524 -3182 -490 -3034
rect -490 -3182 -481 -3034
rect -629 -3410 -620 -3262
rect -620 -3410 -586 -3262
rect -586 -3410 -577 -3262
rect -629 -3422 -577 -3410
rect -341 -3034 -289 -3022
rect -341 -3182 -332 -3034
rect -332 -3182 -298 -3034
rect -298 -3182 -289 -3034
rect -437 -3410 -428 -3262
rect -428 -3410 -394 -3262
rect -394 -3410 -385 -3262
rect -437 -3422 -385 -3410
rect -149 -3034 -97 -3022
rect -149 -3182 -140 -3034
rect -140 -3182 -106 -3034
rect -106 -3182 -97 -3034
rect -245 -3410 -236 -3262
rect -236 -3410 -202 -3262
rect -202 -3410 -193 -3262
rect -245 -3422 -193 -3410
rect 43 -3034 95 -3022
rect 43 -3182 52 -3034
rect 52 -3182 86 -3034
rect 86 -3182 95 -3034
rect -53 -3410 -44 -3262
rect -44 -3410 -10 -3262
rect -10 -3410 -1 -3262
rect -53 -3422 -1 -3410
rect 235 -3034 287 -3022
rect 235 -3182 244 -3034
rect 244 -3182 278 -3034
rect 278 -3182 287 -3034
rect 139 -3410 148 -3262
rect 148 -3410 182 -3262
rect 182 -3410 191 -3262
rect 139 -3422 191 -3410
rect 427 -3034 479 -3022
rect 427 -3182 436 -3034
rect 436 -3182 470 -3034
rect 470 -3182 479 -3034
rect 331 -3410 340 -3262
rect 340 -3410 374 -3262
rect 374 -3410 383 -3262
rect 331 -3422 383 -3410
rect 619 -3034 671 -3022
rect 619 -3182 628 -3034
rect 628 -3182 662 -3034
rect 662 -3182 671 -3034
rect 523 -3410 532 -3262
rect 532 -3410 566 -3262
rect 566 -3410 575 -3262
rect 523 -3422 575 -3410
rect 811 -3034 863 -3022
rect 811 -3182 820 -3034
rect 820 -3182 854 -3034
rect 854 -3182 863 -3034
rect 715 -3410 724 -3262
rect 724 -3410 758 -3262
rect 758 -3410 767 -3262
rect 715 -3422 767 -3410
rect 1003 -3034 1055 -3022
rect 1003 -3182 1012 -3034
rect 1012 -3182 1046 -3034
rect 1046 -3182 1055 -3034
rect 907 -3410 916 -3262
rect 916 -3410 950 -3262
rect 950 -3410 959 -3262
rect 907 -3422 959 -3410
rect 1195 -3034 1247 -3022
rect 1195 -3182 1204 -3034
rect 1204 -3182 1238 -3034
rect 1238 -3182 1247 -3034
rect 1099 -3410 1108 -3262
rect 1108 -3410 1142 -3262
rect 1142 -3410 1151 -3262
rect 1099 -3422 1151 -3410
rect -1205 -3652 -1153 -3640
rect -1205 -3800 -1196 -3652
rect -1196 -3800 -1162 -3652
rect -1162 -3800 -1153 -3652
rect -1380 -4120 -1270 -4020
rect -1013 -3652 -961 -3640
rect -1013 -3800 -1004 -3652
rect -1004 -3800 -970 -3652
rect -970 -3800 -961 -3652
rect -1109 -4028 -1100 -3880
rect -1100 -4028 -1066 -3880
rect -1066 -4028 -1057 -3880
rect -1109 -4040 -1057 -4028
rect -821 -3652 -769 -3640
rect -821 -3800 -812 -3652
rect -812 -3800 -778 -3652
rect -778 -3800 -769 -3652
rect -917 -4028 -908 -3880
rect -908 -4028 -874 -3880
rect -874 -4028 -865 -3880
rect -917 -4040 -865 -4028
rect -629 -3652 -577 -3640
rect -629 -3800 -620 -3652
rect -620 -3800 -586 -3652
rect -586 -3800 -577 -3652
rect -725 -4028 -716 -3880
rect -716 -4028 -682 -3880
rect -682 -4028 -673 -3880
rect -725 -4040 -673 -4028
rect -437 -3652 -385 -3640
rect -437 -3800 -428 -3652
rect -428 -3800 -394 -3652
rect -394 -3800 -385 -3652
rect -533 -4028 -524 -3880
rect -524 -4028 -490 -3880
rect -490 -4028 -481 -3880
rect -533 -4040 -481 -4028
rect -245 -3652 -193 -3640
rect -245 -3800 -236 -3652
rect -236 -3800 -202 -3652
rect -202 -3800 -193 -3652
rect -341 -4028 -332 -3880
rect -332 -4028 -298 -3880
rect -298 -4028 -289 -3880
rect -341 -4040 -289 -4028
rect -53 -3652 -1 -3640
rect -53 -3800 -44 -3652
rect -44 -3800 -10 -3652
rect -10 -3800 -1 -3652
rect -149 -4028 -140 -3880
rect -140 -4028 -106 -3880
rect -106 -4028 -97 -3880
rect -149 -4040 -97 -4028
rect 139 -3652 191 -3640
rect 139 -3800 148 -3652
rect 148 -3800 182 -3652
rect 182 -3800 191 -3652
rect 43 -4028 52 -3880
rect 52 -4028 86 -3880
rect 86 -4028 95 -3880
rect 43 -4040 95 -4028
rect 331 -3652 383 -3640
rect 331 -3800 340 -3652
rect 340 -3800 374 -3652
rect 374 -3800 383 -3652
rect 235 -4028 244 -3880
rect 244 -4028 278 -3880
rect 278 -4028 287 -3880
rect 235 -4040 287 -4028
rect 523 -3652 575 -3640
rect 523 -3800 532 -3652
rect 532 -3800 566 -3652
rect 566 -3800 575 -3652
rect 427 -4028 436 -3880
rect 436 -4028 470 -3880
rect 470 -4028 479 -3880
rect 427 -4040 479 -4028
rect 715 -3652 767 -3640
rect 715 -3800 724 -3652
rect 724 -3800 758 -3652
rect 758 -3800 767 -3652
rect 619 -4028 628 -3880
rect 628 -4028 662 -3880
rect 662 -4028 671 -3880
rect 619 -4040 671 -4028
rect 907 -3652 959 -3640
rect 907 -3800 916 -3652
rect 916 -3800 950 -3652
rect 950 -3800 959 -3652
rect 811 -4028 820 -3880
rect 820 -4028 854 -3880
rect 854 -4028 863 -3880
rect 811 -4040 863 -4028
rect 1099 -3652 1151 -3640
rect 1099 -3800 1108 -3652
rect 1108 -3800 1142 -3652
rect 1142 -3800 1151 -3652
rect 1003 -4028 1012 -3880
rect 1012 -4028 1046 -3880
rect 1046 -4028 1055 -3880
rect 1003 -4040 1055 -4028
rect 1195 -4028 1204 -3880
rect 1204 -4028 1238 -3880
rect 1238 -4028 1247 -3880
rect 1195 -4040 1247 -4028
rect -1087 -4537 -1035 -4525
rect -1087 -4685 -1078 -4537
rect -1078 -4685 -1044 -4537
rect -1044 -4685 -1035 -4537
rect -1185 -4913 -1176 -4765
rect -1176 -4913 -1142 -4765
rect -1142 -4913 -1133 -4765
rect -1185 -4925 -1133 -4913
rect -891 -4537 -839 -4525
rect -891 -4685 -882 -4537
rect -882 -4685 -848 -4537
rect -848 -4685 -839 -4537
rect -989 -4913 -980 -4765
rect -980 -4913 -946 -4765
rect -946 -4913 -937 -4765
rect -989 -4925 -937 -4913
rect -695 -4537 -643 -4525
rect -695 -4685 -686 -4537
rect -686 -4685 -652 -4537
rect -652 -4685 -643 -4537
rect -793 -4913 -784 -4765
rect -784 -4913 -750 -4765
rect -750 -4913 -741 -4765
rect -793 -4925 -741 -4913
rect -499 -4537 -447 -4525
rect -499 -4685 -490 -4537
rect -490 -4685 -456 -4537
rect -456 -4685 -447 -4537
rect -597 -4913 -588 -4765
rect -588 -4913 -554 -4765
rect -554 -4913 -545 -4765
rect -597 -4925 -545 -4913
rect -303 -4537 -251 -4525
rect -303 -4685 -294 -4537
rect -294 -4685 -260 -4537
rect -260 -4685 -251 -4537
rect -401 -4913 -392 -4765
rect -392 -4913 -358 -4765
rect -358 -4913 -349 -4765
rect -401 -4925 -349 -4913
rect -107 -4537 -55 -4525
rect -107 -4685 -98 -4537
rect -98 -4685 -64 -4537
rect -64 -4685 -55 -4537
rect -205 -4913 -196 -4765
rect -196 -4913 -162 -4765
rect -162 -4913 -153 -4765
rect -205 -4925 -153 -4913
rect 89 -4537 141 -4525
rect 89 -4685 98 -4537
rect 98 -4685 132 -4537
rect 132 -4685 141 -4537
rect -9 -4913 0 -4765
rect 0 -4913 34 -4765
rect 34 -4913 43 -4765
rect -9 -4925 43 -4913
rect 285 -4537 337 -4525
rect 285 -4685 294 -4537
rect 294 -4685 328 -4537
rect 328 -4685 337 -4537
rect 187 -4913 196 -4765
rect 196 -4913 230 -4765
rect 230 -4913 239 -4765
rect 187 -4925 239 -4913
rect 711 -4537 763 -4525
rect 711 -4685 720 -4537
rect 720 -4685 754 -4537
rect 754 -4685 763 -4537
rect 613 -4913 622 -4765
rect 622 -4913 656 -4765
rect 656 -4913 665 -4765
rect 613 -4925 665 -4913
rect 907 -4537 959 -4525
rect 907 -4685 916 -4537
rect 916 -4685 950 -4537
rect 950 -4685 959 -4537
rect 809 -4913 818 -4765
rect 818 -4913 852 -4765
rect 852 -4913 861 -4765
rect 809 -4925 861 -4913
rect 1103 -4537 1155 -4525
rect 1103 -4685 1112 -4537
rect 1112 -4685 1146 -4537
rect 1146 -4685 1155 -4537
rect 1005 -4913 1014 -4765
rect 1014 -4913 1048 -4765
rect 1048 -4913 1057 -4765
rect 1005 -4925 1057 -4913
rect 1299 -4537 1351 -4525
rect 1299 -4685 1308 -4537
rect 1308 -4685 1342 -4537
rect 1342 -4685 1351 -4537
rect 1201 -4913 1210 -4765
rect 1210 -4913 1244 -4765
rect 1244 -4913 1253 -4765
rect 1201 -4925 1253 -4913
rect 1495 -4537 1547 -4525
rect 1495 -4685 1504 -4537
rect 1504 -4685 1538 -4537
rect 1538 -4685 1547 -4537
rect 1397 -4913 1406 -4765
rect 1406 -4913 1440 -4765
rect 1440 -4913 1449 -4765
rect 1397 -4925 1449 -4913
rect 1691 -4537 1743 -4525
rect 1691 -4685 1700 -4537
rect 1700 -4685 1734 -4537
rect 1734 -4685 1743 -4537
rect 1593 -4913 1602 -4765
rect 1602 -4913 1636 -4765
rect 1636 -4913 1645 -4765
rect 1593 -4925 1645 -4913
rect 1887 -4537 1939 -4525
rect 1887 -4685 1896 -4537
rect 1896 -4685 1930 -4537
rect 1930 -4685 1939 -4537
rect 1789 -4913 1798 -4765
rect 1798 -4913 1832 -4765
rect 1832 -4913 1841 -4765
rect 1789 -4925 1841 -4913
rect 2083 -4537 2135 -4525
rect 2083 -4685 2092 -4537
rect 2092 -4685 2126 -4537
rect 2126 -4685 2135 -4537
rect 1985 -4913 1994 -4765
rect 1994 -4913 2028 -4765
rect 2028 -4913 2037 -4765
rect 1985 -4925 2037 -4913
rect -1185 -5173 -1133 -5161
rect -1185 -5321 -1176 -5173
rect -1176 -5321 -1142 -5173
rect -1142 -5321 -1133 -5173
rect -989 -5173 -937 -5161
rect -989 -5321 -980 -5173
rect -980 -5321 -946 -5173
rect -946 -5321 -937 -5173
rect -1087 -5549 -1078 -5401
rect -1078 -5549 -1044 -5401
rect -1044 -5549 -1035 -5401
rect -1087 -5561 -1035 -5549
rect -793 -5173 -741 -5161
rect -793 -5321 -784 -5173
rect -784 -5321 -750 -5173
rect -750 -5321 -741 -5173
rect -891 -5549 -882 -5401
rect -882 -5549 -848 -5401
rect -848 -5549 -839 -5401
rect -891 -5561 -839 -5549
rect -597 -5173 -545 -5161
rect -597 -5321 -588 -5173
rect -588 -5321 -554 -5173
rect -554 -5321 -545 -5173
rect -695 -5549 -686 -5401
rect -686 -5549 -652 -5401
rect -652 -5549 -643 -5401
rect -695 -5561 -643 -5549
rect -401 -5173 -349 -5161
rect -401 -5321 -392 -5173
rect -392 -5321 -358 -5173
rect -358 -5321 -349 -5173
rect -499 -5549 -490 -5401
rect -490 -5549 -456 -5401
rect -456 -5549 -447 -5401
rect -499 -5561 -447 -5549
rect -205 -5173 -153 -5161
rect -205 -5321 -196 -5173
rect -196 -5321 -162 -5173
rect -162 -5321 -153 -5173
rect -303 -5549 -294 -5401
rect -294 -5549 -260 -5401
rect -260 -5549 -251 -5401
rect -303 -5561 -251 -5549
rect -9 -5173 43 -5161
rect -9 -5321 0 -5173
rect 0 -5321 34 -5173
rect 34 -5321 43 -5173
rect -107 -5549 -98 -5401
rect -98 -5549 -64 -5401
rect -64 -5549 -55 -5401
rect -107 -5561 -55 -5549
rect 187 -5173 239 -5161
rect 187 -5321 196 -5173
rect 196 -5321 230 -5173
rect 230 -5321 239 -5173
rect 89 -5549 98 -5401
rect 98 -5549 132 -5401
rect 132 -5549 141 -5401
rect 89 -5561 141 -5549
rect 285 -5549 294 -5401
rect 294 -5549 328 -5401
rect 328 -5549 337 -5401
rect 285 -5561 337 -5549
rect 613 -5173 665 -5161
rect 613 -5321 622 -5173
rect 622 -5321 656 -5173
rect 656 -5321 665 -5173
rect 809 -5173 861 -5161
rect 809 -5321 818 -5173
rect 818 -5321 852 -5173
rect 852 -5321 861 -5173
rect 711 -5549 720 -5401
rect 720 -5549 754 -5401
rect 754 -5549 763 -5401
rect 711 -5561 763 -5549
rect 1005 -5173 1057 -5161
rect 1005 -5321 1014 -5173
rect 1014 -5321 1048 -5173
rect 1048 -5321 1057 -5173
rect 907 -5549 916 -5401
rect 916 -5549 950 -5401
rect 950 -5549 959 -5401
rect 907 -5561 959 -5549
rect 1201 -5173 1253 -5161
rect 1201 -5321 1210 -5173
rect 1210 -5321 1244 -5173
rect 1244 -5321 1253 -5173
rect 1103 -5549 1112 -5401
rect 1112 -5549 1146 -5401
rect 1146 -5549 1155 -5401
rect 1103 -5561 1155 -5549
rect 1397 -5173 1449 -5161
rect 1397 -5321 1406 -5173
rect 1406 -5321 1440 -5173
rect 1440 -5321 1449 -5173
rect 1299 -5549 1308 -5401
rect 1308 -5549 1342 -5401
rect 1342 -5549 1351 -5401
rect 1299 -5561 1351 -5549
rect 1593 -5173 1645 -5161
rect 1593 -5321 1602 -5173
rect 1602 -5321 1636 -5173
rect 1636 -5321 1645 -5173
rect 1495 -5549 1504 -5401
rect 1504 -5549 1538 -5401
rect 1538 -5549 1547 -5401
rect 1495 -5561 1547 -5549
rect 1789 -5173 1841 -5161
rect 1789 -5321 1798 -5173
rect 1798 -5321 1832 -5173
rect 1832 -5321 1841 -5173
rect 1691 -5549 1700 -5401
rect 1700 -5549 1734 -5401
rect 1734 -5549 1743 -5401
rect 1691 -5561 1743 -5549
rect 1985 -5173 2037 -5161
rect 1985 -5321 1994 -5173
rect 1994 -5321 2028 -5173
rect 2028 -5321 2037 -5173
rect 1887 -5549 1896 -5401
rect 1896 -5549 1930 -5401
rect 1930 -5549 1939 -5401
rect 1887 -5561 1939 -5549
rect 2083 -5549 2092 -5401
rect 2092 -5549 2126 -5401
rect 2126 -5549 2135 -5401
rect 2083 -5561 2135 -5549
rect 2214 -5560 2344 -5000
rect 2573 -5189 2625 -5177
rect 2573 -5337 2582 -5189
rect 2582 -5337 2616 -5189
rect 2616 -5337 2625 -5189
rect 2415 -5565 2424 -5417
rect 2424 -5565 2458 -5417
rect 2458 -5565 2467 -5417
rect 2415 -5577 2467 -5565
rect 2889 -5189 2941 -5177
rect 2889 -5337 2898 -5189
rect 2898 -5337 2932 -5189
rect 2932 -5337 2941 -5189
rect 2731 -5565 2740 -5417
rect 2740 -5565 2774 -5417
rect 2774 -5565 2783 -5417
rect 2731 -5577 2783 -5565
rect 3205 -5189 3257 -5177
rect 3205 -5337 3214 -5189
rect 3214 -5337 3248 -5189
rect 3248 -5337 3257 -5189
rect 3047 -5565 3056 -5417
rect 3056 -5565 3090 -5417
rect 3090 -5565 3099 -5417
rect 3047 -5577 3099 -5565
rect 3521 -5189 3573 -5177
rect 3521 -5337 3530 -5189
rect 3530 -5337 3564 -5189
rect 3564 -5337 3573 -5189
rect 3363 -5565 3372 -5417
rect 3372 -5565 3406 -5417
rect 3406 -5565 3415 -5417
rect 3363 -5577 3415 -5565
rect 3837 -5189 3889 -5177
rect 3837 -5337 3846 -5189
rect 3846 -5337 3880 -5189
rect 3880 -5337 3889 -5189
rect 3679 -5565 3688 -5417
rect 3688 -5565 3722 -5417
rect 3722 -5565 3731 -5417
rect 3679 -5577 3731 -5565
rect 3995 -5565 4004 -5417
rect 4004 -5565 4038 -5417
rect 4038 -5565 4047 -5417
rect 3995 -5577 4047 -5565
rect 4190 -5200 4290 -5080
rect -1087 -6004 -1035 -5992
rect -1087 -6152 -1078 -6004
rect -1078 -6152 -1044 -6004
rect -1044 -6152 -1035 -6004
rect -1185 -6380 -1176 -6232
rect -1176 -6380 -1142 -6232
rect -1142 -6380 -1133 -6232
rect -1185 -6392 -1133 -6380
rect -891 -6004 -839 -5992
rect -891 -6152 -882 -6004
rect -882 -6152 -848 -6004
rect -848 -6152 -839 -6004
rect -989 -6380 -980 -6232
rect -980 -6380 -946 -6232
rect -946 -6380 -937 -6232
rect -989 -6392 -937 -6380
rect -695 -6004 -643 -5992
rect -695 -6152 -686 -6004
rect -686 -6152 -652 -6004
rect -652 -6152 -643 -6004
rect -793 -6380 -784 -6232
rect -784 -6380 -750 -6232
rect -750 -6380 -741 -6232
rect -793 -6392 -741 -6380
rect -499 -6004 -447 -5992
rect -499 -6152 -490 -6004
rect -490 -6152 -456 -6004
rect -456 -6152 -447 -6004
rect -597 -6380 -588 -6232
rect -588 -6380 -554 -6232
rect -554 -6380 -545 -6232
rect -597 -6392 -545 -6380
rect -303 -6004 -251 -5992
rect -303 -6152 -294 -6004
rect -294 -6152 -260 -6004
rect -260 -6152 -251 -6004
rect -401 -6380 -392 -6232
rect -392 -6380 -358 -6232
rect -358 -6380 -349 -6232
rect -401 -6392 -349 -6380
rect -107 -6004 -55 -5992
rect -107 -6152 -98 -6004
rect -98 -6152 -64 -6004
rect -64 -6152 -55 -6004
rect -205 -6380 -196 -6232
rect -196 -6380 -162 -6232
rect -162 -6380 -153 -6232
rect -205 -6392 -153 -6380
rect 89 -6004 141 -5992
rect 89 -6152 98 -6004
rect 98 -6152 132 -6004
rect 132 -6152 141 -6004
rect -9 -6380 0 -6232
rect 0 -6380 34 -6232
rect 34 -6380 43 -6232
rect -9 -6392 43 -6380
rect 285 -6004 337 -5992
rect 285 -6152 294 -6004
rect 294 -6152 328 -6004
rect 328 -6152 337 -6004
rect 187 -6380 196 -6232
rect 196 -6380 230 -6232
rect 230 -6380 239 -6232
rect 187 -6392 239 -6380
rect 481 -6004 533 -5992
rect 481 -6152 490 -6004
rect 490 -6152 524 -6004
rect 524 -6152 533 -6004
rect 383 -6380 392 -6232
rect 392 -6380 426 -6232
rect 426 -6380 435 -6232
rect 383 -6392 435 -6380
rect 677 -6004 729 -5992
rect 677 -6152 686 -6004
rect 686 -6152 720 -6004
rect 720 -6152 729 -6004
rect 579 -6380 588 -6232
rect 588 -6380 622 -6232
rect 622 -6380 631 -6232
rect 579 -6392 631 -6380
rect 873 -6004 925 -5992
rect 873 -6152 882 -6004
rect 882 -6152 916 -6004
rect 916 -6152 925 -6004
rect 775 -6380 784 -6232
rect 784 -6380 818 -6232
rect 818 -6380 827 -6232
rect 775 -6392 827 -6380
rect 1069 -6004 1121 -5992
rect 1069 -6152 1078 -6004
rect 1078 -6152 1112 -6004
rect 1112 -6152 1121 -6004
rect 971 -6380 980 -6232
rect 980 -6380 1014 -6232
rect 1014 -6380 1023 -6232
rect 971 -6392 1023 -6380
rect 1265 -6004 1317 -5992
rect 1265 -6152 1274 -6004
rect 1274 -6152 1308 -6004
rect 1308 -6152 1317 -6004
rect 1167 -6380 1176 -6232
rect 1176 -6380 1210 -6232
rect 1210 -6380 1219 -6232
rect 1167 -6392 1219 -6380
rect 2164 -6410 2414 -6220
rect -1185 -6622 -1133 -6610
rect -1185 -6770 -1176 -6622
rect -1176 -6770 -1142 -6622
rect -1142 -6770 -1133 -6622
rect -989 -6622 -937 -6610
rect -989 -6770 -980 -6622
rect -980 -6770 -946 -6622
rect -946 -6770 -937 -6622
rect -1087 -6998 -1078 -6850
rect -1078 -6998 -1044 -6850
rect -1044 -6998 -1035 -6850
rect -1087 -7010 -1035 -6998
rect -793 -6622 -741 -6610
rect -793 -6770 -784 -6622
rect -784 -6770 -750 -6622
rect -750 -6770 -741 -6622
rect -891 -6998 -882 -6850
rect -882 -6998 -848 -6850
rect -848 -6998 -839 -6850
rect -891 -7010 -839 -6998
rect -597 -6622 -545 -6610
rect -597 -6770 -588 -6622
rect -588 -6770 -554 -6622
rect -554 -6770 -545 -6622
rect -695 -6998 -686 -6850
rect -686 -6998 -652 -6850
rect -652 -6998 -643 -6850
rect -695 -7010 -643 -6998
rect -401 -6622 -349 -6610
rect -401 -6770 -392 -6622
rect -392 -6770 -358 -6622
rect -358 -6770 -349 -6622
rect -499 -6998 -490 -6850
rect -490 -6998 -456 -6850
rect -456 -6998 -447 -6850
rect -499 -7010 -447 -6998
rect -205 -6622 -153 -6610
rect -205 -6770 -196 -6622
rect -196 -6770 -162 -6622
rect -162 -6770 -153 -6622
rect -303 -6998 -294 -6850
rect -294 -6998 -260 -6850
rect -260 -6998 -251 -6850
rect -303 -7010 -251 -6998
rect -9 -6622 43 -6610
rect -9 -6770 0 -6622
rect 0 -6770 34 -6622
rect 34 -6770 43 -6622
rect -107 -6998 -98 -6850
rect -98 -6998 -64 -6850
rect -64 -6998 -55 -6850
rect -107 -7010 -55 -6998
rect 187 -6622 239 -6610
rect 187 -6770 196 -6622
rect 196 -6770 230 -6622
rect 230 -6770 239 -6622
rect 89 -6998 98 -6850
rect 98 -6998 132 -6850
rect 132 -6998 141 -6850
rect 89 -7010 141 -6998
rect 383 -6622 435 -6610
rect 383 -6770 392 -6622
rect 392 -6770 426 -6622
rect 426 -6770 435 -6622
rect 285 -6998 294 -6850
rect 294 -6998 328 -6850
rect 328 -6998 337 -6850
rect 285 -7010 337 -6998
rect 579 -6622 631 -6610
rect 579 -6770 588 -6622
rect 588 -6770 622 -6622
rect 622 -6770 631 -6622
rect 481 -6998 490 -6850
rect 490 -6998 524 -6850
rect 524 -6998 533 -6850
rect 481 -7010 533 -6998
rect 775 -6622 827 -6610
rect 775 -6770 784 -6622
rect 784 -6770 818 -6622
rect 818 -6770 827 -6622
rect 677 -6998 686 -6850
rect 686 -6998 720 -6850
rect 720 -6998 729 -6850
rect 677 -7010 729 -6998
rect 971 -6622 1023 -6610
rect 971 -6770 980 -6622
rect 980 -6770 1014 -6622
rect 1014 -6770 1023 -6622
rect 873 -6998 882 -6850
rect 882 -6998 916 -6850
rect 916 -6998 925 -6850
rect 873 -7010 925 -6998
rect 1167 -6622 1219 -6610
rect 1167 -6770 1176 -6622
rect 1176 -6770 1210 -6622
rect 1210 -6770 1219 -6622
rect 1069 -6998 1078 -6850
rect 1078 -6998 1112 -6850
rect 1112 -6998 1121 -6850
rect 1069 -7010 1121 -6998
rect 2475 -6324 2527 -6312
rect 2475 -6472 2484 -6324
rect 2484 -6472 2518 -6324
rect 2518 -6472 2527 -6324
rect 2671 -6324 2723 -6312
rect 2671 -6472 2680 -6324
rect 2680 -6472 2714 -6324
rect 2714 -6472 2723 -6324
rect 2573 -6700 2582 -6552
rect 2582 -6700 2616 -6552
rect 2616 -6700 2625 -6552
rect 2573 -6712 2625 -6700
rect 2867 -6324 2919 -6312
rect 2867 -6472 2876 -6324
rect 2876 -6472 2910 -6324
rect 2910 -6472 2919 -6324
rect 2769 -6700 2778 -6552
rect 2778 -6700 2812 -6552
rect 2812 -6700 2821 -6552
rect 2769 -6712 2821 -6700
rect 3063 -6324 3115 -6312
rect 3063 -6472 3072 -6324
rect 3072 -6472 3106 -6324
rect 3106 -6472 3115 -6324
rect 2965 -6700 2974 -6552
rect 2974 -6700 3008 -6552
rect 3008 -6700 3017 -6552
rect 2965 -6712 3017 -6700
rect 3259 -6324 3311 -6312
rect 3259 -6472 3268 -6324
rect 3268 -6472 3302 -6324
rect 3302 -6472 3311 -6324
rect 3161 -6700 3170 -6552
rect 3170 -6700 3204 -6552
rect 3204 -6700 3213 -6552
rect 3161 -6712 3213 -6700
rect 3455 -6324 3507 -6312
rect 3455 -6472 3464 -6324
rect 3464 -6472 3498 -6324
rect 3498 -6472 3507 -6324
rect 3357 -6700 3366 -6552
rect 3366 -6700 3400 -6552
rect 3400 -6700 3409 -6552
rect 3357 -6712 3409 -6700
rect 3651 -6324 3703 -6312
rect 3651 -6472 3660 -6324
rect 3660 -6472 3694 -6324
rect 3694 -6472 3703 -6324
rect 3553 -6700 3562 -6552
rect 3562 -6700 3596 -6552
rect 3596 -6700 3605 -6552
rect 3553 -6712 3605 -6700
rect 3847 -6324 3899 -6312
rect 3847 -6472 3856 -6324
rect 3856 -6472 3890 -6324
rect 3890 -6472 3899 -6324
rect 3749 -6700 3758 -6552
rect 3758 -6700 3792 -6552
rect 3792 -6700 3801 -6552
rect 3749 -6712 3801 -6700
rect 3945 -6700 3954 -6552
rect 3954 -6700 3988 -6552
rect 3988 -6700 3997 -6552
rect 3945 -6712 3997 -6700
rect 1265 -6998 1274 -6850
rect 1274 -6998 1308 -6850
rect 1308 -6998 1317 -6850
rect 1265 -7010 1317 -6998
rect 1454 -6910 1684 -6750
rect 2204 -6910 2284 -6750
rect -1087 -7448 -1035 -7436
rect -1087 -7596 -1078 -7448
rect -1078 -7596 -1044 -7448
rect -1044 -7596 -1035 -7448
rect -1185 -7824 -1176 -7676
rect -1176 -7824 -1142 -7676
rect -1142 -7824 -1133 -7676
rect -1185 -7836 -1133 -7824
rect -891 -7448 -839 -7436
rect -891 -7596 -882 -7448
rect -882 -7596 -848 -7448
rect -848 -7596 -839 -7448
rect -989 -7824 -980 -7676
rect -980 -7824 -946 -7676
rect -946 -7824 -937 -7676
rect -989 -7836 -937 -7824
rect -695 -7448 -643 -7436
rect -695 -7596 -686 -7448
rect -686 -7596 -652 -7448
rect -652 -7596 -643 -7448
rect -793 -7824 -784 -7676
rect -784 -7824 -750 -7676
rect -750 -7824 -741 -7676
rect -793 -7836 -741 -7824
rect -499 -7448 -447 -7436
rect -499 -7596 -490 -7448
rect -490 -7596 -456 -7448
rect -456 -7596 -447 -7448
rect -597 -7824 -588 -7676
rect -588 -7824 -554 -7676
rect -554 -7824 -545 -7676
rect -597 -7836 -545 -7824
rect -303 -7448 -251 -7436
rect -303 -7596 -294 -7448
rect -294 -7596 -260 -7448
rect -260 -7596 -251 -7448
rect -401 -7824 -392 -7676
rect -392 -7824 -358 -7676
rect -358 -7824 -349 -7676
rect -401 -7836 -349 -7824
rect -107 -7448 -55 -7436
rect -107 -7596 -98 -7448
rect -98 -7596 -64 -7448
rect -64 -7596 -55 -7448
rect -205 -7824 -196 -7676
rect -196 -7824 -162 -7676
rect -162 -7824 -153 -7676
rect -205 -7836 -153 -7824
rect 89 -7448 141 -7436
rect 89 -7596 98 -7448
rect 98 -7596 132 -7448
rect 132 -7596 141 -7448
rect -9 -7824 0 -7676
rect 0 -7824 34 -7676
rect 34 -7824 43 -7676
rect -9 -7836 43 -7824
rect 285 -7448 337 -7436
rect 285 -7596 294 -7448
rect 294 -7596 328 -7448
rect 328 -7596 337 -7448
rect 187 -7824 196 -7676
rect 196 -7824 230 -7676
rect 230 -7824 239 -7676
rect 187 -7836 239 -7824
rect 481 -7448 533 -7436
rect 481 -7596 490 -7448
rect 490 -7596 524 -7448
rect 524 -7596 533 -7448
rect 383 -7824 392 -7676
rect 392 -7824 426 -7676
rect 426 -7824 435 -7676
rect 383 -7836 435 -7824
rect 677 -7448 729 -7436
rect 677 -7596 686 -7448
rect 686 -7596 720 -7448
rect 720 -7596 729 -7448
rect 579 -7824 588 -7676
rect 588 -7824 622 -7676
rect 622 -7824 631 -7676
rect 579 -7836 631 -7824
rect 873 -7448 925 -7436
rect 873 -7596 882 -7448
rect 882 -7596 916 -7448
rect 916 -7596 925 -7448
rect 775 -7824 784 -7676
rect 784 -7824 818 -7676
rect 818 -7824 827 -7676
rect 775 -7836 827 -7824
rect 1069 -7448 1121 -7436
rect 1069 -7596 1078 -7448
rect 1078 -7596 1112 -7448
rect 1112 -7596 1121 -7448
rect 971 -7824 980 -7676
rect 980 -7824 1014 -7676
rect 1014 -7824 1023 -7676
rect 971 -7836 1023 -7824
rect 1265 -7448 1317 -7436
rect 1265 -7596 1274 -7448
rect 1274 -7596 1308 -7448
rect 1308 -7596 1317 -7448
rect 1167 -7824 1176 -7676
rect 1176 -7824 1210 -7676
rect 1210 -7824 1219 -7676
rect 1167 -7836 1219 -7824
rect 2573 -6942 2625 -6930
rect 2573 -7090 2582 -6942
rect 2582 -7090 2616 -6942
rect 2616 -7090 2625 -6942
rect 2475 -7318 2484 -7170
rect 2484 -7318 2518 -7170
rect 2518 -7318 2527 -7170
rect 2475 -7330 2527 -7318
rect 2769 -6942 2821 -6930
rect 2769 -7090 2778 -6942
rect 2778 -7090 2812 -6942
rect 2812 -7090 2821 -6942
rect 2671 -7318 2680 -7170
rect 2680 -7318 2714 -7170
rect 2714 -7318 2723 -7170
rect 2671 -7330 2723 -7318
rect 2965 -6942 3017 -6930
rect 2965 -7090 2974 -6942
rect 2974 -7090 3008 -6942
rect 3008 -7090 3017 -6942
rect 2867 -7318 2876 -7170
rect 2876 -7318 2910 -7170
rect 2910 -7318 2919 -7170
rect 2867 -7330 2919 -7318
rect 3161 -6942 3213 -6930
rect 3161 -7090 3170 -6942
rect 3170 -7090 3204 -6942
rect 3204 -7090 3213 -6942
rect 3063 -7318 3072 -7170
rect 3072 -7318 3106 -7170
rect 3106 -7318 3115 -7170
rect 3063 -7330 3115 -7318
rect 3357 -6942 3409 -6930
rect 3357 -7090 3366 -6942
rect 3366 -7090 3400 -6942
rect 3400 -7090 3409 -6942
rect 3259 -7318 3268 -7170
rect 3268 -7318 3302 -7170
rect 3302 -7318 3311 -7170
rect 3259 -7330 3311 -7318
rect 3553 -6942 3605 -6930
rect 3553 -7090 3562 -6942
rect 3562 -7090 3596 -6942
rect 3596 -7090 3605 -6942
rect 3455 -7318 3464 -7170
rect 3464 -7318 3498 -7170
rect 3498 -7318 3507 -7170
rect 3455 -7330 3507 -7318
rect 3749 -6942 3801 -6930
rect 3749 -7090 3758 -6942
rect 3758 -7090 3792 -6942
rect 3792 -7090 3801 -6942
rect 3651 -7318 3660 -7170
rect 3660 -7318 3694 -7170
rect 3694 -7318 3703 -7170
rect 3651 -7330 3703 -7318
rect 3945 -6942 3997 -6930
rect 3945 -7090 3954 -6942
rect 3954 -7090 3988 -6942
rect 3988 -7090 3997 -6942
rect 4054 -6940 4174 -6730
rect 3847 -7318 3856 -7170
rect 3856 -7318 3890 -7170
rect 3890 -7318 3899 -7170
rect 3847 -7330 3899 -7318
rect -1185 -8066 -1133 -8054
rect -1185 -8214 -1176 -8066
rect -1176 -8214 -1142 -8066
rect -1142 -8214 -1133 -8066
rect -989 -8066 -937 -8054
rect -989 -8214 -980 -8066
rect -980 -8214 -946 -8066
rect -946 -8214 -937 -8066
rect -1087 -8442 -1078 -8294
rect -1078 -8442 -1044 -8294
rect -1044 -8442 -1035 -8294
rect -1087 -8454 -1035 -8442
rect -793 -8066 -741 -8054
rect -793 -8214 -784 -8066
rect -784 -8214 -750 -8066
rect -750 -8214 -741 -8066
rect -891 -8442 -882 -8294
rect -882 -8442 -848 -8294
rect -848 -8442 -839 -8294
rect -891 -8454 -839 -8442
rect -597 -8066 -545 -8054
rect -597 -8214 -588 -8066
rect -588 -8214 -554 -8066
rect -554 -8214 -545 -8066
rect -695 -8442 -686 -8294
rect -686 -8442 -652 -8294
rect -652 -8442 -643 -8294
rect -695 -8454 -643 -8442
rect -401 -8066 -349 -8054
rect -401 -8214 -392 -8066
rect -392 -8214 -358 -8066
rect -358 -8214 -349 -8066
rect -499 -8442 -490 -8294
rect -490 -8442 -456 -8294
rect -456 -8442 -447 -8294
rect -499 -8454 -447 -8442
rect -205 -8066 -153 -8054
rect -205 -8214 -196 -8066
rect -196 -8214 -162 -8066
rect -162 -8214 -153 -8066
rect -303 -8442 -294 -8294
rect -294 -8442 -260 -8294
rect -260 -8442 -251 -8294
rect -303 -8454 -251 -8442
rect -9 -8066 43 -8054
rect -9 -8214 0 -8066
rect 0 -8214 34 -8066
rect 34 -8214 43 -8066
rect -107 -8442 -98 -8294
rect -98 -8442 -64 -8294
rect -64 -8442 -55 -8294
rect -107 -8454 -55 -8442
rect 187 -8066 239 -8054
rect 187 -8214 196 -8066
rect 196 -8214 230 -8066
rect 230 -8214 239 -8066
rect 89 -8442 98 -8294
rect 98 -8442 132 -8294
rect 132 -8442 141 -8294
rect 89 -8454 141 -8442
rect 383 -8066 435 -8054
rect 383 -8214 392 -8066
rect 392 -8214 426 -8066
rect 426 -8214 435 -8066
rect 285 -8442 294 -8294
rect 294 -8442 328 -8294
rect 328 -8442 337 -8294
rect 285 -8454 337 -8442
rect 579 -8066 631 -8054
rect 579 -8214 588 -8066
rect 588 -8214 622 -8066
rect 622 -8214 631 -8066
rect 481 -8442 490 -8294
rect 490 -8442 524 -8294
rect 524 -8442 533 -8294
rect 481 -8454 533 -8442
rect 775 -8066 827 -8054
rect 775 -8214 784 -8066
rect 784 -8214 818 -8066
rect 818 -8214 827 -8066
rect 677 -8442 686 -8294
rect 686 -8442 720 -8294
rect 720 -8442 729 -8294
rect 677 -8454 729 -8442
rect 971 -8066 1023 -8054
rect 971 -8214 980 -8066
rect 980 -8214 1014 -8066
rect 1014 -8214 1023 -8066
rect 873 -8442 882 -8294
rect 882 -8442 916 -8294
rect 916 -8442 925 -8294
rect 873 -8454 925 -8442
rect 1167 -8066 1219 -8054
rect 1167 -8214 1176 -8066
rect 1176 -8214 1210 -8066
rect 1210 -8214 1219 -8066
rect 1069 -8442 1078 -8294
rect 1078 -8442 1112 -8294
rect 1112 -8442 1121 -8294
rect 1069 -8454 1121 -8442
rect 1265 -8442 1274 -8294
rect 1274 -8442 1308 -8294
rect 1308 -8442 1317 -8294
rect 1265 -8454 1317 -8442
rect 1701 -8102 1753 -8090
rect 1701 -8250 1710 -8102
rect 1710 -8250 1744 -8102
rect 1744 -8250 1753 -8102
rect 1605 -8478 1614 -8330
rect 1614 -8478 1648 -8330
rect 1648 -8478 1657 -8330
rect 1605 -8490 1657 -8478
rect 1893 -8102 1945 -8090
rect 1893 -8250 1902 -8102
rect 1902 -8250 1936 -8102
rect 1936 -8250 1945 -8102
rect 1797 -8478 1806 -8330
rect 1806 -8478 1840 -8330
rect 1840 -8478 1849 -8330
rect 1797 -8490 1849 -8478
rect 2085 -8102 2137 -8090
rect 2085 -8250 2094 -8102
rect 2094 -8250 2128 -8102
rect 2128 -8250 2137 -8102
rect 1989 -8478 1998 -8330
rect 1998 -8478 2032 -8330
rect 2032 -8478 2041 -8330
rect 1989 -8490 2041 -8478
rect 2277 -8102 2329 -8090
rect 2277 -8250 2286 -8102
rect 2286 -8250 2320 -8102
rect 2320 -8250 2329 -8102
rect 2181 -8478 2190 -8330
rect 2190 -8478 2224 -8330
rect 2224 -8478 2233 -8330
rect 2181 -8490 2233 -8478
rect 2469 -8102 2521 -8090
rect 2469 -8250 2478 -8102
rect 2478 -8250 2512 -8102
rect 2512 -8250 2521 -8102
rect 2373 -8478 2382 -8330
rect 2382 -8478 2416 -8330
rect 2416 -8478 2425 -8330
rect 2373 -8490 2425 -8478
rect 2661 -8102 2713 -8090
rect 2661 -8250 2670 -8102
rect 2670 -8250 2704 -8102
rect 2704 -8250 2713 -8102
rect 2565 -8478 2574 -8330
rect 2574 -8478 2608 -8330
rect 2608 -8478 2617 -8330
rect 2565 -8490 2617 -8478
rect 2850 -8140 3020 -7990
rect 2757 -8478 2766 -8330
rect 2766 -8478 2800 -8330
rect 2800 -8478 2809 -8330
rect 2757 -8490 2809 -8478
rect 3597 -8102 3649 -8090
rect 3597 -8250 3606 -8102
rect 3606 -8250 3640 -8102
rect 3640 -8250 3649 -8102
rect 3501 -8478 3510 -8330
rect 3510 -8478 3544 -8330
rect 3544 -8478 3553 -8330
rect 3501 -8490 3553 -8478
rect 3789 -8102 3841 -8090
rect 3789 -8250 3798 -8102
rect 3798 -8250 3832 -8102
rect 3832 -8250 3841 -8102
rect 3693 -8478 3702 -8330
rect 3702 -8478 3736 -8330
rect 3736 -8478 3745 -8330
rect 3693 -8490 3745 -8478
rect 3981 -8102 4033 -8090
rect 3981 -8250 3990 -8102
rect 3990 -8250 4024 -8102
rect 4024 -8250 4033 -8102
rect 3885 -8478 3894 -8330
rect 3894 -8478 3928 -8330
rect 3928 -8478 3937 -8330
rect 3885 -8490 3937 -8478
rect 4173 -8102 4225 -8090
rect 4173 -8250 4182 -8102
rect 4182 -8250 4216 -8102
rect 4216 -8250 4225 -8102
rect 4077 -8478 4086 -8330
rect 4086 -8478 4120 -8330
rect 4120 -8478 4129 -8330
rect 4077 -8490 4129 -8478
rect 4365 -8102 4417 -8090
rect 4365 -8250 4374 -8102
rect 4374 -8250 4408 -8102
rect 4408 -8250 4417 -8102
rect 4269 -8478 4278 -8330
rect 4278 -8478 4312 -8330
rect 4312 -8478 4321 -8330
rect 4269 -8490 4321 -8478
rect 4557 -8102 4609 -8090
rect 4557 -8250 4566 -8102
rect 4566 -8250 4600 -8102
rect 4600 -8250 4609 -8102
rect 4461 -8478 4470 -8330
rect 4470 -8478 4504 -8330
rect 4504 -8478 4513 -8330
rect 4461 -8490 4513 -8478
rect 4653 -8478 4662 -8330
rect 4662 -8478 4696 -8330
rect 4696 -8478 4705 -8330
rect 4653 -8490 4705 -8478
rect -1380 -8850 -1270 -8760
rect -1109 -8868 -1057 -8856
rect -1109 -9016 -1100 -8868
rect -1100 -9016 -1066 -8868
rect -1066 -9016 -1057 -8868
rect -1205 -9244 -1196 -9096
rect -1196 -9244 -1162 -9096
rect -1162 -9244 -1153 -9096
rect -1205 -9256 -1153 -9244
rect -917 -8868 -865 -8856
rect -917 -9016 -908 -8868
rect -908 -9016 -874 -8868
rect -874 -9016 -865 -8868
rect -1013 -9244 -1004 -9096
rect -1004 -9244 -970 -9096
rect -970 -9244 -961 -9096
rect -1013 -9256 -961 -9244
rect -725 -8868 -673 -8856
rect -725 -9016 -716 -8868
rect -716 -9016 -682 -8868
rect -682 -9016 -673 -8868
rect -821 -9244 -812 -9096
rect -812 -9244 -778 -9096
rect -778 -9244 -769 -9096
rect -821 -9256 -769 -9244
rect -533 -8868 -481 -8856
rect -533 -9016 -524 -8868
rect -524 -9016 -490 -8868
rect -490 -9016 -481 -8868
rect -629 -9244 -620 -9096
rect -620 -9244 -586 -9096
rect -586 -9244 -577 -9096
rect -629 -9256 -577 -9244
rect -341 -8868 -289 -8856
rect -341 -9016 -332 -8868
rect -332 -9016 -298 -8868
rect -298 -9016 -289 -8868
rect -437 -9244 -428 -9096
rect -428 -9244 -394 -9096
rect -394 -9244 -385 -9096
rect -437 -9256 -385 -9244
rect -149 -8868 -97 -8856
rect -149 -9016 -140 -8868
rect -140 -9016 -106 -8868
rect -106 -9016 -97 -8868
rect -245 -9244 -236 -9096
rect -236 -9244 -202 -9096
rect -202 -9244 -193 -9096
rect -245 -9256 -193 -9244
rect 43 -8868 95 -8856
rect 43 -9016 52 -8868
rect 52 -9016 86 -8868
rect 86 -9016 95 -8868
rect -53 -9244 -44 -9096
rect -44 -9244 -10 -9096
rect -10 -9244 -1 -9096
rect -53 -9256 -1 -9244
rect 235 -8868 287 -8856
rect 235 -9016 244 -8868
rect 244 -9016 278 -8868
rect 278 -9016 287 -8868
rect 139 -9244 148 -9096
rect 148 -9244 182 -9096
rect 182 -9244 191 -9096
rect 139 -9256 191 -9244
rect 427 -8868 479 -8856
rect 427 -9016 436 -8868
rect 436 -9016 470 -8868
rect 470 -9016 479 -8868
rect 331 -9244 340 -9096
rect 340 -9244 374 -9096
rect 374 -9244 383 -9096
rect 331 -9256 383 -9244
rect 619 -8868 671 -8856
rect 619 -9016 628 -8868
rect 628 -9016 662 -8868
rect 662 -9016 671 -8868
rect 523 -9244 532 -9096
rect 532 -9244 566 -9096
rect 566 -9244 575 -9096
rect 523 -9256 575 -9244
rect 811 -8868 863 -8856
rect 811 -9016 820 -8868
rect 820 -9016 854 -8868
rect 854 -9016 863 -8868
rect 715 -9244 724 -9096
rect 724 -9244 758 -9096
rect 758 -9244 767 -9096
rect 715 -9256 767 -9244
rect 1003 -8868 1055 -8856
rect 1003 -9016 1012 -8868
rect 1012 -9016 1046 -8868
rect 1046 -9016 1055 -8868
rect 907 -9244 916 -9096
rect 916 -9244 950 -9096
rect 950 -9244 959 -9096
rect 907 -9256 959 -9244
rect 1195 -8868 1247 -8856
rect 1195 -9016 1204 -8868
rect 1204 -9016 1238 -8868
rect 1238 -9016 1247 -8868
rect 1099 -9244 1108 -9096
rect 1108 -9244 1142 -9096
rect 1142 -9244 1151 -9096
rect 1099 -9256 1151 -9244
rect 1344 -9320 1474 -9140
rect 1863 -8922 1915 -8910
rect 1863 -9070 1872 -8922
rect 1872 -9070 1906 -8922
rect 1906 -9070 1915 -8922
rect 1605 -9298 1614 -9150
rect 1614 -9298 1648 -9150
rect 1648 -9298 1657 -9150
rect 1605 -9310 1657 -9298
rect 2379 -8922 2431 -8910
rect 2379 -9070 2388 -8922
rect 2388 -9070 2422 -8922
rect 2422 -9070 2431 -8922
rect 2121 -9298 2130 -9150
rect 2130 -9298 2164 -9150
rect 2164 -9298 2173 -9150
rect 2121 -9310 2173 -9298
rect 2895 -8922 2947 -8910
rect 2895 -9070 2904 -8922
rect 2904 -9070 2938 -8922
rect 2938 -9070 2947 -8922
rect 2637 -9298 2646 -9150
rect 2646 -9298 2680 -9150
rect 2680 -9298 2689 -9150
rect 2637 -9310 2689 -9298
rect 3759 -8922 3811 -8910
rect 3759 -9070 3768 -8922
rect 3768 -9070 3802 -8922
rect 3802 -9070 3811 -8922
rect 3153 -9298 3162 -9150
rect 3162 -9298 3196 -9150
rect 3196 -9298 3205 -9150
rect 3153 -9310 3205 -9298
rect 3501 -9298 3510 -9150
rect 3510 -9298 3544 -9150
rect 3544 -9298 3553 -9150
rect 3501 -9310 3553 -9298
rect 4275 -8922 4327 -8910
rect 4275 -9070 4284 -8922
rect 4284 -9070 4318 -8922
rect 4318 -9070 4327 -8922
rect 4017 -9298 4026 -9150
rect 4026 -9298 4060 -9150
rect 4060 -9298 4069 -9150
rect 4017 -9310 4069 -9298
rect 4791 -8922 4843 -8910
rect 4791 -9070 4800 -8922
rect 4800 -9070 4834 -8922
rect 4834 -9070 4843 -8922
rect 4533 -9298 4542 -9150
rect 4542 -9298 4576 -9150
rect 4576 -9298 4585 -9150
rect 4533 -9310 4585 -9298
rect 5440 -8922 5500 -8910
rect 5440 -9090 5460 -8922
rect 5460 -9090 5494 -8922
rect 5494 -9090 5500 -8922
rect 5049 -9298 5058 -9150
rect 5058 -9298 5092 -9150
rect 5092 -9298 5101 -9150
rect 5049 -9310 5101 -9298
rect 5640 -8922 5700 -8910
rect 5640 -9090 5652 -8922
rect 5652 -9090 5686 -8922
rect 5686 -9090 5700 -8922
rect 5540 -9298 5556 -9150
rect 5556 -9298 5590 -9150
rect 5590 -9298 5600 -9150
rect 5540 -9310 5600 -9298
rect 5830 -8922 5890 -8910
rect 5830 -9090 5844 -8922
rect 5844 -9090 5878 -8922
rect 5878 -9090 5890 -8922
rect 5740 -9298 5748 -9150
rect 5748 -9298 5782 -9150
rect 5782 -9298 5800 -9150
rect 5740 -9310 5800 -9298
rect 5930 -9298 5940 -9150
rect 5940 -9298 5974 -9150
rect 5974 -9298 5990 -9150
rect 5930 -9310 5990 -9298
rect 6060 -9410 6130 -9300
rect -1205 -9486 -1153 -9474
rect -1205 -9634 -1196 -9486
rect -1196 -9634 -1162 -9486
rect -1162 -9634 -1153 -9486
rect -1013 -9486 -961 -9474
rect -1013 -9634 -1004 -9486
rect -1004 -9634 -970 -9486
rect -970 -9634 -961 -9486
rect -1109 -9862 -1100 -9714
rect -1100 -9862 -1066 -9714
rect -1066 -9862 -1057 -9714
rect -1109 -9874 -1057 -9862
rect -821 -9486 -769 -9474
rect -821 -9634 -812 -9486
rect -812 -9634 -778 -9486
rect -778 -9634 -769 -9486
rect -917 -9862 -908 -9714
rect -908 -9862 -874 -9714
rect -874 -9862 -865 -9714
rect -917 -9874 -865 -9862
rect -629 -9486 -577 -9474
rect -629 -9634 -620 -9486
rect -620 -9634 -586 -9486
rect -586 -9634 -577 -9486
rect -725 -9862 -716 -9714
rect -716 -9862 -682 -9714
rect -682 -9862 -673 -9714
rect -725 -9874 -673 -9862
rect -437 -9486 -385 -9474
rect -437 -9634 -428 -9486
rect -428 -9634 -394 -9486
rect -394 -9634 -385 -9486
rect -533 -9862 -524 -9714
rect -524 -9862 -490 -9714
rect -490 -9862 -481 -9714
rect -533 -9874 -481 -9862
rect -245 -9486 -193 -9474
rect -245 -9634 -236 -9486
rect -236 -9634 -202 -9486
rect -202 -9634 -193 -9486
rect -341 -9862 -332 -9714
rect -332 -9862 -298 -9714
rect -298 -9862 -289 -9714
rect -341 -9874 -289 -9862
rect -53 -9486 -1 -9474
rect -53 -9634 -44 -9486
rect -44 -9634 -10 -9486
rect -10 -9634 -1 -9486
rect -149 -9862 -140 -9714
rect -140 -9862 -106 -9714
rect -106 -9862 -97 -9714
rect -149 -9874 -97 -9862
rect 139 -9486 191 -9474
rect 139 -9634 148 -9486
rect 148 -9634 182 -9486
rect 182 -9634 191 -9486
rect 43 -9862 52 -9714
rect 52 -9862 86 -9714
rect 86 -9862 95 -9714
rect 43 -9874 95 -9862
rect 331 -9486 383 -9474
rect 331 -9634 340 -9486
rect 340 -9634 374 -9486
rect 374 -9634 383 -9486
rect 235 -9862 244 -9714
rect 244 -9862 278 -9714
rect 278 -9862 287 -9714
rect 235 -9874 287 -9862
rect 523 -9486 575 -9474
rect 523 -9634 532 -9486
rect 532 -9634 566 -9486
rect 566 -9634 575 -9486
rect 427 -9862 436 -9714
rect 436 -9862 470 -9714
rect 470 -9862 479 -9714
rect 427 -9874 479 -9862
rect 715 -9486 767 -9474
rect 715 -9634 724 -9486
rect 724 -9634 758 -9486
rect 758 -9634 767 -9486
rect 619 -9862 628 -9714
rect 628 -9862 662 -9714
rect 662 -9862 671 -9714
rect 619 -9874 671 -9862
rect 907 -9486 959 -9474
rect 907 -9634 916 -9486
rect 916 -9634 950 -9486
rect 950 -9634 959 -9486
rect 811 -9862 820 -9714
rect 820 -9862 854 -9714
rect 854 -9862 863 -9714
rect 811 -9874 863 -9862
rect 1099 -9486 1151 -9474
rect 1099 -9634 1108 -9486
rect 1108 -9634 1142 -9486
rect 1142 -9634 1151 -9486
rect 1003 -9862 1012 -9714
rect 1012 -9862 1046 -9714
rect 1046 -9862 1055 -9714
rect 1003 -9874 1055 -9862
rect 1195 -9862 1204 -9714
rect 1204 -9862 1238 -9714
rect 1238 -9862 1247 -9714
rect 1195 -9874 1247 -9862
rect -1109 -10104 -1057 -10092
rect -1109 -10252 -1100 -10104
rect -1100 -10252 -1066 -10104
rect -1066 -10252 -1057 -10104
rect -1205 -10480 -1196 -10332
rect -1196 -10480 -1162 -10332
rect -1162 -10480 -1153 -10332
rect -1205 -10492 -1153 -10480
rect -917 -10104 -865 -10092
rect -917 -10252 -908 -10104
rect -908 -10252 -874 -10104
rect -874 -10252 -865 -10104
rect -1013 -10480 -1004 -10332
rect -1004 -10480 -970 -10332
rect -970 -10480 -961 -10332
rect -1013 -10492 -961 -10480
rect -725 -10104 -673 -10092
rect -725 -10252 -716 -10104
rect -716 -10252 -682 -10104
rect -682 -10252 -673 -10104
rect -821 -10480 -812 -10332
rect -812 -10480 -778 -10332
rect -778 -10480 -769 -10332
rect -821 -10492 -769 -10480
rect -533 -10104 -481 -10092
rect -533 -10252 -524 -10104
rect -524 -10252 -490 -10104
rect -490 -10252 -481 -10104
rect -629 -10480 -620 -10332
rect -620 -10480 -586 -10332
rect -586 -10480 -577 -10332
rect -629 -10492 -577 -10480
rect -341 -10104 -289 -10092
rect -341 -10252 -332 -10104
rect -332 -10252 -298 -10104
rect -298 -10252 -289 -10104
rect -437 -10480 -428 -10332
rect -428 -10480 -394 -10332
rect -394 -10480 -385 -10332
rect -437 -10492 -385 -10480
rect -149 -10104 -97 -10092
rect -149 -10252 -140 -10104
rect -140 -10252 -106 -10104
rect -106 -10252 -97 -10104
rect -245 -10480 -236 -10332
rect -236 -10480 -202 -10332
rect -202 -10480 -193 -10332
rect -245 -10492 -193 -10480
rect 43 -10104 95 -10092
rect 43 -10252 52 -10104
rect 52 -10252 86 -10104
rect 86 -10252 95 -10104
rect -53 -10480 -44 -10332
rect -44 -10480 -10 -10332
rect -10 -10480 -1 -10332
rect -53 -10492 -1 -10480
rect 235 -10104 287 -10092
rect 235 -10252 244 -10104
rect 244 -10252 278 -10104
rect 278 -10252 287 -10104
rect 139 -10480 148 -10332
rect 148 -10480 182 -10332
rect 182 -10480 191 -10332
rect 139 -10492 191 -10480
rect 427 -10104 479 -10092
rect 427 -10252 436 -10104
rect 436 -10252 470 -10104
rect 470 -10252 479 -10104
rect 331 -10480 340 -10332
rect 340 -10480 374 -10332
rect 374 -10480 383 -10332
rect 331 -10492 383 -10480
rect 619 -10104 671 -10092
rect 619 -10252 628 -10104
rect 628 -10252 662 -10104
rect 662 -10252 671 -10104
rect 523 -10480 532 -10332
rect 532 -10480 566 -10332
rect 566 -10480 575 -10332
rect 523 -10492 575 -10480
rect 811 -10104 863 -10092
rect 811 -10252 820 -10104
rect 820 -10252 854 -10104
rect 854 -10252 863 -10104
rect 715 -10480 724 -10332
rect 724 -10480 758 -10332
rect 758 -10480 767 -10332
rect 715 -10492 767 -10480
rect 1003 -10104 1055 -10092
rect 1003 -10252 1012 -10104
rect 1012 -10252 1046 -10104
rect 1046 -10252 1055 -10104
rect 907 -10480 916 -10332
rect 916 -10480 950 -10332
rect 950 -10480 959 -10332
rect 907 -10492 959 -10480
rect 1195 -10104 1247 -10092
rect 1195 -10252 1204 -10104
rect 1204 -10252 1238 -10104
rect 1238 -10252 1247 -10104
rect 1099 -10480 1108 -10332
rect 1108 -10480 1142 -10332
rect 1142 -10480 1151 -10332
rect 1099 -10492 1151 -10480
rect -1205 -10722 -1153 -10710
rect -1205 -10870 -1196 -10722
rect -1196 -10870 -1162 -10722
rect -1162 -10870 -1153 -10722
rect -1013 -10722 -961 -10710
rect -1013 -10870 -1004 -10722
rect -1004 -10870 -970 -10722
rect -970 -10870 -961 -10722
rect -1109 -11098 -1100 -10950
rect -1100 -11098 -1066 -10950
rect -1066 -11098 -1057 -10950
rect -1109 -11110 -1057 -11098
rect -821 -10722 -769 -10710
rect -821 -10870 -812 -10722
rect -812 -10870 -778 -10722
rect -778 -10870 -769 -10722
rect -917 -11098 -908 -10950
rect -908 -11098 -874 -10950
rect -874 -11098 -865 -10950
rect -917 -11110 -865 -11098
rect -629 -10722 -577 -10710
rect -629 -10870 -620 -10722
rect -620 -10870 -586 -10722
rect -586 -10870 -577 -10722
rect -725 -11098 -716 -10950
rect -716 -11098 -682 -10950
rect -682 -11098 -673 -10950
rect -725 -11110 -673 -11098
rect -437 -10722 -385 -10710
rect -437 -10870 -428 -10722
rect -428 -10870 -394 -10722
rect -394 -10870 -385 -10722
rect -533 -11098 -524 -10950
rect -524 -11098 -490 -10950
rect -490 -11098 -481 -10950
rect -533 -11110 -481 -11098
rect -245 -10722 -193 -10710
rect -245 -10870 -236 -10722
rect -236 -10870 -202 -10722
rect -202 -10870 -193 -10722
rect -341 -11098 -332 -10950
rect -332 -11098 -298 -10950
rect -298 -11098 -289 -10950
rect -341 -11110 -289 -11098
rect -53 -10722 -1 -10710
rect -53 -10870 -44 -10722
rect -44 -10870 -10 -10722
rect -10 -10870 -1 -10722
rect -149 -11098 -140 -10950
rect -140 -11098 -106 -10950
rect -106 -11098 -97 -10950
rect -149 -11110 -97 -11098
rect 139 -10722 191 -10710
rect 139 -10870 148 -10722
rect 148 -10870 182 -10722
rect 182 -10870 191 -10722
rect 43 -11098 52 -10950
rect 52 -11098 86 -10950
rect 86 -11098 95 -10950
rect 43 -11110 95 -11098
rect 331 -10722 383 -10710
rect 331 -10870 340 -10722
rect 340 -10870 374 -10722
rect 374 -10870 383 -10722
rect 235 -11098 244 -10950
rect 244 -11098 278 -10950
rect 278 -11098 287 -10950
rect 235 -11110 287 -11098
rect 523 -10722 575 -10710
rect 523 -10870 532 -10722
rect 532 -10870 566 -10722
rect 566 -10870 575 -10722
rect 427 -11098 436 -10950
rect 436 -11098 470 -10950
rect 470 -11098 479 -10950
rect 427 -11110 479 -11098
rect 715 -10722 767 -10710
rect 715 -10870 724 -10722
rect 724 -10870 758 -10722
rect 758 -10870 767 -10722
rect 619 -11098 628 -10950
rect 628 -11098 662 -10950
rect 662 -11098 671 -10950
rect 619 -11110 671 -11098
rect 907 -10722 959 -10710
rect 907 -10870 916 -10722
rect 916 -10870 950 -10722
rect 950 -10870 959 -10722
rect 811 -11098 820 -10950
rect 820 -11098 854 -10950
rect 854 -11098 863 -10950
rect 811 -11110 863 -11098
rect 1099 -10722 1151 -10710
rect 1099 -10870 1108 -10722
rect 1108 -10870 1142 -10722
rect 1142 -10870 1151 -10722
rect 1003 -11098 1012 -10950
rect 1012 -11098 1046 -10950
rect 1046 -11098 1055 -10950
rect 1003 -11110 1055 -11098
rect 1195 -11098 1204 -10950
rect 1204 -11098 1238 -10950
rect 1238 -11098 1247 -10950
rect 1195 -11110 1247 -11098
rect 6390 -10070 6460 -9960
rect 6620 -10223 6670 -10200
rect 6620 -10299 6622 -10223
rect 6622 -10299 6670 -10223
rect 6620 -10320 6670 -10299
rect 6670 -10320 6760 -10200
<< metal2 >>
rect -1087 2550 -1035 2555
rect -891 2550 -839 2555
rect -695 2550 -643 2555
rect -499 2550 -447 2555
rect -303 2550 -251 2555
rect -107 2550 -55 2555
rect 89 2550 141 2555
rect 285 2550 337 2555
rect 711 2550 763 2555
rect 907 2550 959 2555
rect 1103 2550 1155 2555
rect 1299 2550 1351 2555
rect 1495 2550 1547 2555
rect 1691 2550 1743 2555
rect 1887 2550 1939 2555
rect 2083 2550 2135 2555
rect -1096 2545 2304 2550
rect -1096 2385 -1087 2545
rect -1035 2385 -891 2545
rect -839 2385 -695 2545
rect -643 2385 -499 2545
rect -447 2385 -303 2545
rect -251 2385 -107 2545
rect -55 2385 89 2545
rect 141 2385 285 2545
rect 337 2530 711 2545
rect 337 2390 354 2530
rect 594 2390 711 2530
rect 337 2385 711 2390
rect 763 2385 907 2545
rect 959 2385 1103 2545
rect 1155 2385 1299 2545
rect 1351 2385 1495 2545
rect 1547 2385 1691 2545
rect 1743 2385 1887 2545
rect 1939 2385 2083 2545
rect 2135 2385 2304 2545
rect -1096 2380 2304 2385
rect -1087 2375 -1035 2380
rect -891 2375 -839 2380
rect -695 2375 -643 2380
rect -499 2375 -447 2380
rect -303 2375 -251 2380
rect -107 2375 -55 2380
rect 89 2375 141 2380
rect 285 2375 337 2380
rect 711 2375 763 2380
rect 907 2375 959 2380
rect 1103 2375 1155 2380
rect 1299 2375 1351 2380
rect 1495 2375 1547 2380
rect 1691 2375 1743 2380
rect 1887 2375 1939 2380
rect 2054 2370 2304 2380
rect -1185 2310 -1133 2315
rect -989 2310 -937 2315
rect -793 2310 -741 2315
rect -597 2310 -545 2315
rect -401 2310 -349 2315
rect -205 2310 -153 2315
rect -9 2310 43 2315
rect 187 2310 239 2315
rect 613 2310 665 2315
rect 809 2310 861 2315
rect 1005 2310 1057 2315
rect 1201 2310 1253 2315
rect 1397 2310 1449 2315
rect 1593 2310 1645 2315
rect 1789 2310 1841 2315
rect 1985 2310 2037 2315
rect -1196 2305 2044 2310
rect -1196 2145 -1185 2305
rect -1133 2145 -989 2305
rect -937 2145 -793 2305
rect -741 2145 -597 2305
rect -545 2145 -401 2305
rect -349 2145 -205 2305
rect -153 2145 -9 2305
rect 43 2145 187 2305
rect 239 2145 613 2305
rect 665 2145 809 2305
rect 861 2300 1005 2305
rect 1057 2300 1201 2305
rect 1253 2300 1397 2305
rect 861 2150 974 2300
rect 1374 2150 1397 2300
rect 861 2145 1005 2150
rect 1057 2145 1201 2150
rect 1253 2145 1397 2150
rect 1449 2145 1593 2305
rect 1645 2145 1789 2305
rect 1841 2145 1985 2305
rect 2037 2145 2044 2305
rect -1196 2140 2044 2145
rect -1185 2135 -1133 2140
rect -989 2135 -937 2140
rect -793 2135 -741 2140
rect -597 2135 -545 2140
rect -401 2135 -349 2140
rect -205 2135 -153 2140
rect -9 2135 43 2140
rect 187 2135 239 2140
rect 613 2135 665 2140
rect 809 2135 861 2140
rect 1005 2135 1057 2140
rect 1201 2135 1253 2140
rect 1397 2135 1449 2140
rect 1593 2135 1645 2140
rect 1789 2135 1841 2140
rect 1985 2135 2037 2140
rect 2164 2090 2304 2370
rect 2164 2070 3894 2090
rect -1185 1910 -1133 1919
rect -989 1910 -937 1919
rect -793 1910 -741 1919
rect -597 1910 -545 1919
rect -401 1910 -349 1919
rect -205 1910 -153 1919
rect -9 1910 43 1919
rect 187 1910 239 1919
rect 613 1910 665 1919
rect 809 1910 861 1919
rect 1005 1910 1057 1919
rect 1201 1910 1253 1919
rect 1397 1910 1449 1919
rect 1593 1910 1645 1919
rect 1789 1910 1841 1919
rect 1985 1910 2037 1919
rect -1196 1909 2044 1910
rect -1196 1749 -1185 1909
rect -1133 1749 -989 1909
rect -937 1749 -793 1909
rect -741 1749 -597 1909
rect -545 1749 -401 1909
rect -349 1749 -205 1909
rect -153 1749 -9 1909
rect 43 1749 187 1909
rect 239 1749 613 1909
rect 665 1749 809 1909
rect 861 1900 1005 1909
rect 1057 1900 1201 1909
rect 1253 1900 1397 1909
rect 861 1750 984 1900
rect 1384 1750 1397 1900
rect 861 1749 1005 1750
rect 1057 1749 1201 1750
rect 1253 1749 1397 1750
rect 1449 1749 1593 1909
rect 1645 1749 1789 1909
rect 1841 1749 1985 1909
rect 2037 1749 2044 1909
rect -1196 1740 2044 1749
rect -1185 1739 -1133 1740
rect -989 1739 -937 1740
rect -793 1739 -741 1740
rect -597 1739 -545 1740
rect -401 1739 -349 1740
rect -205 1739 -153 1740
rect -9 1739 43 1740
rect 187 1739 239 1740
rect 613 1739 665 1740
rect 809 1739 861 1740
rect 1005 1739 1057 1740
rect 1201 1739 1253 1740
rect 1397 1739 1449 1740
rect 1593 1739 1645 1740
rect 1789 1739 1841 1740
rect 1985 1739 2037 1740
rect 2164 1680 2214 2070
rect -1087 1670 -1035 1679
rect -891 1670 -839 1679
rect -695 1670 -643 1679
rect -499 1670 -447 1679
rect -303 1670 -251 1679
rect -107 1670 -55 1679
rect 89 1670 141 1679
rect 285 1670 337 1679
rect 711 1670 763 1679
rect 907 1670 959 1679
rect 1103 1670 1155 1679
rect 1299 1670 1351 1679
rect 1495 1670 1547 1679
rect 1691 1670 1743 1679
rect 1887 1670 1939 1679
rect 2054 1670 2214 1680
rect -1087 1669 2214 1670
rect -1035 1510 -891 1669
rect -1087 1499 -1035 1509
rect -839 1510 -695 1669
rect -891 1499 -839 1509
rect -643 1510 -499 1669
rect -695 1499 -643 1509
rect -447 1510 -303 1669
rect -499 1499 -447 1509
rect -251 1510 -107 1669
rect -303 1499 -251 1509
rect -55 1510 89 1669
rect -107 1499 -55 1509
rect 141 1510 285 1669
rect 89 1499 141 1509
rect 337 1650 711 1669
rect 337 1510 354 1650
rect 594 1510 711 1650
rect 337 1509 614 1510
rect 285 1499 614 1509
rect 763 1510 907 1669
rect 711 1499 763 1509
rect 959 1510 1103 1669
rect 907 1499 959 1509
rect 1155 1510 1299 1669
rect 1103 1499 1155 1509
rect 1351 1510 1495 1669
rect 1299 1499 1351 1509
rect 1547 1510 1691 1669
rect 1495 1499 1547 1509
rect 1743 1510 1887 1669
rect 1691 1499 1743 1509
rect 1939 1510 2083 1669
rect 1887 1499 1939 1509
rect 2135 1510 2214 1669
rect 2344 1893 3894 2070
rect 4660 2000 4740 2010
rect 4660 1920 4740 1930
rect 2344 1733 2573 1893
rect 2625 1733 2889 1893
rect 2941 1733 3205 1893
rect 3257 1733 3521 1893
rect 3573 1733 3837 1893
rect 3889 1733 3894 1893
rect 2344 1730 3894 1733
rect 2573 1723 2625 1730
rect 2889 1723 2941 1730
rect 3205 1723 3257 1730
rect 3521 1723 3573 1730
rect 3837 1723 3889 1730
rect 2834 1670 3274 1680
rect 2415 1660 2467 1663
rect 2731 1660 2783 1663
rect 2083 1499 2135 1509
rect 2214 1500 2344 1510
rect 2414 1653 2834 1660
rect 3363 1660 3415 1663
rect 3679 1660 3731 1663
rect 3995 1660 4047 1663
rect 3274 1653 4054 1660
rect 314 1490 614 1499
rect 2414 1493 2415 1653
rect 2467 1493 2731 1653
rect 2783 1493 2834 1653
rect 3274 1493 3363 1653
rect 3415 1493 3679 1653
rect 3731 1493 3995 1653
rect 4047 1493 4054 1653
rect 2414 1490 2834 1493
rect 3274 1490 4054 1493
rect 2415 1483 2467 1490
rect 2731 1483 2783 1490
rect 2834 1480 3274 1490
rect 3363 1483 3415 1490
rect 3679 1483 3731 1490
rect 3995 1483 4047 1490
rect 524 1088 844 1090
rect -1087 1080 -1035 1088
rect -891 1080 -839 1088
rect -695 1080 -643 1088
rect -499 1080 -447 1088
rect -303 1080 -251 1088
rect -107 1080 -55 1088
rect 89 1080 141 1088
rect 285 1080 337 1088
rect 481 1080 844 1088
rect 873 1080 925 1088
rect 1069 1080 1121 1088
rect 1265 1080 1317 1088
rect -1096 1078 524 1080
rect 844 1078 1324 1080
rect -1096 918 -1087 1078
rect -1035 918 -891 1078
rect -839 918 -695 1078
rect -643 918 -499 1078
rect -447 918 -303 1078
rect -251 918 -107 1078
rect -55 918 89 1078
rect 141 918 285 1078
rect 337 918 481 1078
rect 844 918 873 1078
rect 925 918 1069 1078
rect 1121 918 1265 1078
rect 1317 918 1324 1078
rect -1096 910 524 918
rect 844 910 1324 918
rect -1087 908 -1035 910
rect -891 908 -839 910
rect -695 908 -643 910
rect -499 908 -447 910
rect -303 908 -251 910
rect -107 908 -55 910
rect 89 908 141 910
rect 285 908 337 910
rect 481 908 844 910
rect 873 908 925 910
rect 1069 908 1121 910
rect 1265 908 1317 910
rect 524 900 844 908
rect 2164 850 2414 860
rect -1185 840 -1133 848
rect -989 840 -937 848
rect -793 840 -741 848
rect -597 840 -545 848
rect -401 840 -349 848
rect -205 840 -153 848
rect -9 840 43 848
rect 187 840 239 848
rect 383 840 435 848
rect 579 840 631 848
rect 775 840 827 848
rect 971 840 1023 848
rect 1167 840 1219 848
rect -1186 838 2164 840
rect -1186 678 -1185 838
rect -1133 678 -989 838
rect -937 678 -793 838
rect -741 678 -597 838
rect -545 678 -401 838
rect -349 678 -205 838
rect -153 678 -9 838
rect 43 678 187 838
rect 239 678 383 838
rect 435 678 579 838
rect 631 678 775 838
rect 827 678 971 838
rect 1023 830 1167 838
rect 1219 830 2164 838
rect 1384 680 2164 830
rect 1023 678 1167 680
rect 1219 678 2164 680
rect -1186 670 2164 678
rect -1185 668 -1133 670
rect -989 668 -937 670
rect -793 668 -741 670
rect -597 668 -545 670
rect -401 668 -349 670
rect -205 668 -153 670
rect -9 668 43 670
rect 187 668 239 670
rect 383 668 435 670
rect 579 668 631 670
rect 775 668 827 670
rect 971 668 1023 670
rect 1167 668 1219 670
rect 2834 770 3274 780
rect 2164 650 2414 660
rect 2464 758 2834 770
rect 3274 758 3914 770
rect 2464 598 2475 758
rect 2527 598 2671 758
rect 2723 598 2834 758
rect 3311 598 3455 758
rect 3507 598 3651 758
rect 3703 598 3847 758
rect 3899 598 3914 758
rect 2464 590 2834 598
rect 3274 590 3914 598
rect 2475 588 2527 590
rect 2671 588 2723 590
rect 2834 588 3311 590
rect 3455 588 3507 590
rect 3651 588 3703 590
rect 3847 588 3899 590
rect 2834 580 3274 588
rect 2564 518 4114 530
rect -1186 460 1384 470
rect -1186 300 -1185 460
rect -1133 300 -989 460
rect -937 300 -793 460
rect -741 300 -597 460
rect -545 300 -401 460
rect -349 300 -205 460
rect -153 300 -9 460
rect 43 300 187 460
rect 239 300 383 460
rect 435 300 579 460
rect 631 300 775 460
rect 827 300 971 460
rect 2564 358 2573 518
rect 2625 358 2769 518
rect 2821 358 2965 518
rect 3017 358 3161 518
rect 3213 358 3357 518
rect 3409 358 3553 518
rect 3605 358 3749 518
rect 3801 358 3945 518
rect 3997 358 4114 518
rect 2564 350 4114 358
rect 2573 348 2734 350
rect 2769 348 2821 350
rect 2965 348 3017 350
rect 3161 348 3213 350
rect 3357 348 3409 350
rect 3553 348 3605 350
rect 3749 348 3801 350
rect 1023 300 1167 310
rect 1219 300 1384 310
rect 1454 320 1684 330
rect 2204 320 2284 330
rect 2574 320 2734 348
rect 3924 340 4174 350
rect -1185 290 -1133 300
rect -989 290 -937 300
rect -793 290 -741 300
rect -597 290 -545 300
rect -401 290 -349 300
rect -205 290 -153 300
rect -9 290 43 300
rect 187 290 239 300
rect 383 290 435 300
rect 579 290 631 300
rect 775 290 827 300
rect 971 290 1023 300
rect 1167 290 1219 300
rect -1087 220 -1035 230
rect -891 220 -839 230
rect -695 220 -643 230
rect -499 220 -447 230
rect -303 220 -251 230
rect -107 220 -55 230
rect 89 220 141 230
rect 285 220 337 230
rect 424 220 1317 230
rect -1096 60 -1087 220
rect -1035 60 -891 220
rect -839 60 -695 220
rect -643 60 -499 220
rect -447 60 -303 220
rect -251 60 -107 220
rect -55 60 89 220
rect 141 60 285 220
rect 337 60 481 220
rect 844 60 873 220
rect 925 60 1069 220
rect 1121 60 1265 220
rect 1317 60 1324 220
rect 1684 160 2204 320
rect 2284 160 2734 320
rect 1454 150 1684 160
rect 2204 150 2284 160
rect 2564 150 2734 160
rect 4004 150 4054 340
rect -1096 -366 524 60
rect 844 -366 1324 60
rect 2564 140 4054 150
rect 2564 -20 2573 140
rect 2625 -20 2769 140
rect 2821 -20 2965 140
rect 3017 -20 3161 140
rect 3213 -20 3357 140
rect 3409 -20 3553 140
rect 3605 -20 3749 140
rect 3801 -20 3945 140
rect 3997 130 4054 140
rect 3997 120 4174 130
rect 3997 -20 4114 120
rect 2564 -30 4114 -20
rect 2834 -90 3274 -80
rect 2464 -100 2834 -90
rect 3274 -100 3914 -90
rect 2464 -260 2475 -100
rect 2527 -260 2671 -100
rect 2723 -260 2834 -100
rect 3311 -260 3455 -100
rect 3507 -260 3651 -100
rect 3703 -260 3847 -100
rect 3899 -260 3914 -100
rect 2464 -270 2834 -260
rect 3274 -270 3914 -260
rect 2834 -280 3274 -270
rect -1096 -526 -1087 -366
rect -1035 -526 -891 -366
rect -839 -526 -695 -366
rect -643 -526 -499 -366
rect -447 -526 -303 -366
rect -251 -526 -107 -366
rect -55 -526 89 -366
rect 141 -526 285 -366
rect 337 -526 481 -366
rect 844 -526 873 -366
rect 925 -526 1069 -366
rect 1121 -526 1265 -366
rect 1317 -526 1324 -366
rect -1096 -530 524 -526
rect 844 -530 1324 -526
rect -1087 -536 -1035 -530
rect -891 -536 -839 -530
rect -695 -536 -643 -530
rect -499 -536 -447 -530
rect -303 -536 -251 -530
rect -107 -536 -55 -530
rect 89 -536 141 -530
rect 285 -536 337 -530
rect 434 -536 925 -530
rect 1069 -536 1121 -530
rect 1265 -536 1317 -530
rect 434 -540 924 -536
rect -1185 -600 -1133 -596
rect -989 -600 -937 -596
rect -793 -600 -741 -596
rect -597 -600 -545 -596
rect -401 -600 -349 -596
rect -205 -600 -153 -596
rect -9 -600 43 -596
rect 187 -600 239 -596
rect 383 -600 435 -596
rect 579 -600 631 -596
rect 775 -600 827 -596
rect 971 -600 1023 -596
rect 1167 -600 1219 -596
rect -1196 -606 1384 -600
rect -1196 -766 -1185 -606
rect -1133 -766 -989 -606
rect -937 -766 -793 -606
rect -741 -766 -597 -606
rect -545 -766 -401 -606
rect -349 -766 -205 -606
rect -153 -766 -9 -606
rect 43 -766 187 -606
rect 239 -766 383 -606
rect 435 -766 579 -606
rect 631 -766 775 -606
rect 827 -766 971 -606
rect 1023 -610 1167 -606
rect 1219 -610 1384 -606
rect 1023 -766 1167 -760
rect 1219 -766 1384 -760
rect -1196 -770 1384 -766
rect -1185 -776 -1133 -770
rect -989 -776 -937 -770
rect -793 -776 -741 -770
rect -597 -776 -545 -770
rect -401 -776 -349 -770
rect -205 -776 -153 -770
rect -9 -776 43 -770
rect 187 -776 239 -770
rect 383 -776 435 -770
rect 579 -776 631 -770
rect 775 -776 827 -770
rect 971 -776 1023 -770
rect 1167 -776 1219 -770
rect -1186 -980 1804 -970
rect -1186 -984 984 -980
rect -1186 -1140 -1185 -984
rect -1133 -1140 -989 -984
rect -1185 -1154 -1133 -1144
rect -937 -1140 -793 -984
rect -989 -1154 -937 -1144
rect -741 -1140 -597 -984
rect -793 -1154 -741 -1144
rect -545 -1140 -401 -984
rect -597 -1154 -545 -1144
rect -349 -1140 -205 -984
rect -401 -1154 -349 -1144
rect -153 -1140 -9 -984
rect -205 -1154 -153 -1144
rect 43 -1140 187 -984
rect -9 -1154 43 -1144
rect 239 -1140 383 -984
rect 187 -1154 239 -1144
rect 435 -1140 579 -984
rect 383 -1154 435 -1144
rect 631 -1140 775 -984
rect 579 -1154 631 -1144
rect 827 -1140 971 -984
rect 1384 -1010 1804 -980
rect 1384 -1020 2724 -1010
rect 1384 -1130 1701 -1020
rect 775 -1154 827 -1144
rect 1023 -1140 1167 -1130
rect 971 -1154 1023 -1144
rect 1219 -1140 1701 -1130
rect 1167 -1154 1219 -1144
rect 1694 -1180 1701 -1140
rect 1753 -1180 1893 -1020
rect 1945 -1180 2085 -1020
rect 2137 -1180 2277 -1020
rect 2329 -1180 2469 -1020
rect 2521 -1180 2661 -1020
rect 2713 -1180 2724 -1020
rect 1694 -1190 2724 -1180
rect 524 -1214 844 -1210
rect -1087 -1220 -1035 -1214
rect -891 -1220 -839 -1214
rect -695 -1220 -643 -1214
rect -499 -1220 -447 -1214
rect -303 -1220 -251 -1214
rect -107 -1220 -55 -1214
rect 89 -1220 141 -1214
rect 285 -1220 337 -1214
rect 481 -1220 844 -1214
rect 873 -1220 925 -1214
rect 1069 -1220 1121 -1214
rect 1265 -1220 1317 -1214
rect -1096 -1224 524 -1220
rect 844 -1224 1324 -1220
rect -1096 -1384 -1087 -1224
rect -1035 -1384 -891 -1224
rect -839 -1384 -695 -1224
rect -643 -1384 -499 -1224
rect -447 -1384 -303 -1224
rect -251 -1384 -107 -1224
rect -55 -1384 89 -1224
rect 141 -1384 285 -1224
rect 337 -1384 481 -1224
rect 844 -1384 873 -1224
rect 925 -1384 1069 -1224
rect 1121 -1384 1265 -1224
rect 1317 -1384 1324 -1224
rect -1096 -1390 524 -1384
rect 844 -1390 1324 -1384
rect 1604 -1260 2954 -1250
rect -1087 -1394 -1035 -1390
rect -891 -1394 -839 -1390
rect -695 -1394 -643 -1390
rect -499 -1394 -447 -1390
rect -303 -1394 -251 -1390
rect -107 -1394 -55 -1390
rect 89 -1394 141 -1390
rect 285 -1394 337 -1390
rect 481 -1394 844 -1390
rect 873 -1394 925 -1390
rect 1069 -1394 1121 -1390
rect 1265 -1394 1317 -1390
rect 524 -1400 844 -1394
rect 1604 -1420 1605 -1260
rect 1657 -1420 1797 -1260
rect 1849 -1420 1989 -1260
rect 2041 -1420 2181 -1260
rect 2233 -1420 2373 -1260
rect 2425 -1420 2565 -1260
rect 2617 -1420 2757 -1260
rect 2809 -1420 2954 -1260
rect 1604 -1430 2954 -1420
rect -146 -1770 174 -1760
rect -1109 -1780 -1057 -1776
rect -917 -1780 -865 -1776
rect -725 -1780 -673 -1776
rect -533 -1780 -481 -1776
rect -341 -1780 -289 -1776
rect -149 -1780 -146 -1776
rect -1116 -1786 -146 -1780
rect 235 -1780 287 -1776
rect 427 -1780 479 -1776
rect 619 -1780 671 -1776
rect 811 -1780 863 -1776
rect 1003 -1780 1055 -1776
rect 1195 -1780 1247 -1776
rect 174 -1786 1384 -1780
rect -1116 -1946 -1109 -1786
rect -1057 -1946 -917 -1786
rect -865 -1946 -725 -1786
rect -673 -1946 -533 -1786
rect -481 -1946 -341 -1786
rect -289 -1946 -149 -1786
rect 174 -1946 235 -1786
rect 287 -1946 427 -1786
rect 479 -1946 619 -1786
rect 671 -1946 811 -1786
rect 863 -1946 1003 -1786
rect 1055 -1946 1195 -1786
rect 1247 -1946 1384 -1786
rect 2654 -1810 2954 -1430
rect 3140 -1660 3320 -1650
rect 3140 -1790 3320 -1780
rect -1116 -1950 -146 -1946
rect 174 -1950 1384 -1946
rect -1109 -1956 -1057 -1950
rect -917 -1956 -865 -1950
rect -725 -1956 -673 -1950
rect -533 -1956 -481 -1950
rect -341 -1956 -289 -1950
rect -149 -1956 174 -1950
rect 235 -1956 287 -1950
rect 427 -1956 479 -1950
rect 619 -1956 671 -1950
rect 811 -1956 863 -1950
rect 1003 -1956 1055 -1950
rect 1195 -1956 1384 -1950
rect -146 -1960 174 -1956
rect -1205 -2020 -1153 -2016
rect -1013 -2020 -961 -2016
rect -821 -2020 -769 -2016
rect -629 -2020 -577 -2016
rect -437 -2020 -385 -2016
rect -245 -2020 -193 -2016
rect -53 -2020 -1 -2016
rect 139 -2020 191 -2016
rect 331 -2020 383 -2016
rect 523 -2020 575 -2016
rect 715 -2020 767 -2016
rect 907 -2020 959 -2016
rect 1099 -2020 1151 -2016
rect -1216 -2026 1154 -2020
rect -1216 -2186 -1205 -2026
rect -1153 -2186 -1013 -2026
rect -961 -2186 -821 -2026
rect -769 -2186 -629 -2026
rect -577 -2186 -437 -2026
rect -385 -2186 -245 -2026
rect -193 -2186 -53 -2026
rect -1 -2186 139 -2026
rect 191 -2186 331 -2026
rect 383 -2186 523 -2026
rect 575 -2030 715 -2026
rect 767 -2030 907 -2026
rect 844 -2186 907 -2030
rect 959 -2186 1099 -2026
rect 1151 -2186 1154 -2026
rect -1216 -2404 524 -2186
rect 844 -2404 1154 -2186
rect -1216 -2564 -1205 -2404
rect -1153 -2564 -1013 -2404
rect -961 -2564 -821 -2404
rect -769 -2564 -629 -2404
rect -577 -2564 -437 -2404
rect -385 -2564 -245 -2404
rect -193 -2564 -53 -2404
rect -1 -2564 139 -2404
rect 191 -2564 331 -2404
rect 383 -2564 523 -2404
rect 844 -2564 907 -2404
rect 959 -2564 1099 -2404
rect 1151 -2564 1154 -2404
rect -1216 -2570 524 -2564
rect 844 -2570 1154 -2564
rect 1244 -2060 1384 -1956
rect 1844 -1840 2954 -1810
rect 1844 -2000 1863 -1840
rect 1915 -2000 2379 -1840
rect 2431 -2000 2895 -1840
rect 2947 -2000 2954 -1840
rect 1844 -2010 2954 -2000
rect 1244 -2070 1474 -2060
rect 1244 -2150 1344 -2070
rect 1474 -2080 3214 -2070
rect 1474 -2150 1605 -2080
rect 1244 -2420 1260 -2150
rect 1530 -2240 1605 -2150
rect 1657 -2240 2121 -2080
rect 2173 -2240 2637 -2080
rect 2689 -2240 3153 -2080
rect 3205 -2240 3214 -2080
rect 1530 -2250 3214 -2240
rect 1244 -2430 1530 -2420
rect -1205 -2574 -1153 -2570
rect -1013 -2574 -961 -2570
rect -821 -2574 -769 -2570
rect -629 -2574 -577 -2570
rect -437 -2574 -385 -2570
rect -245 -2574 -193 -2570
rect -53 -2574 -1 -2570
rect 139 -2574 191 -2570
rect 331 -2574 383 -2570
rect 523 -2574 844 -2570
rect 907 -2574 959 -2570
rect 1099 -2574 1151 -2570
rect 524 -2580 844 -2574
rect 1244 -2634 1384 -2430
rect -1109 -2640 -1057 -2634
rect -917 -2640 -865 -2634
rect -725 -2640 -673 -2634
rect -533 -2640 -481 -2634
rect -341 -2640 -289 -2634
rect -149 -2640 -97 -2634
rect 43 -2640 95 -2634
rect 235 -2640 287 -2634
rect 427 -2640 479 -2634
rect 619 -2640 671 -2634
rect 811 -2640 863 -2634
rect 1003 -2640 1055 -2634
rect 1195 -2640 1384 -2634
rect -1116 -2644 1384 -2640
rect -1116 -2804 -1109 -2644
rect -1057 -2804 -917 -2644
rect -865 -2804 -725 -2644
rect -673 -2804 -533 -2644
rect -481 -2804 -341 -2644
rect -289 -2804 -149 -2644
rect -97 -2650 43 -2644
rect 95 -2650 235 -2644
rect 174 -2804 235 -2650
rect 287 -2804 427 -2644
rect 479 -2804 619 -2644
rect 671 -2804 811 -2644
rect 863 -2804 1003 -2644
rect 1055 -2804 1195 -2644
rect 1247 -2804 1384 -2644
rect -1116 -3022 -146 -2804
rect 174 -3022 1384 -2804
rect -1116 -3182 -1109 -3022
rect -1057 -3182 -917 -3022
rect -865 -3182 -725 -3022
rect -673 -3182 -533 -3022
rect -481 -3182 -341 -3022
rect -289 -3182 -149 -3022
rect 174 -3182 235 -3022
rect 287 -3182 427 -3022
rect 479 -3182 619 -3022
rect 671 -3182 811 -3022
rect 863 -3182 1003 -3022
rect 1055 -3182 1195 -3022
rect 1247 -3182 1384 -3022
rect -1116 -3190 -146 -3182
rect 174 -3190 1384 -3182
rect -1109 -3192 -1057 -3190
rect -917 -3192 -865 -3190
rect -725 -3192 -673 -3190
rect -533 -3192 -481 -3190
rect -341 -3192 -289 -3190
rect -149 -3192 174 -3190
rect 235 -3192 287 -3190
rect 427 -3192 479 -3190
rect 619 -3192 671 -3190
rect 811 -3192 863 -3190
rect 1003 -3192 1055 -3190
rect 1195 -3192 1384 -3190
rect -146 -3200 174 -3192
rect -1226 -3260 1164 -3250
rect -1226 -3262 524 -3260
rect 844 -3262 1164 -3260
rect -1226 -3422 -1205 -3262
rect -1153 -3422 -1013 -3262
rect -961 -3422 -821 -3262
rect -769 -3422 -629 -3262
rect -577 -3422 -437 -3262
rect -385 -3422 -245 -3262
rect -193 -3422 -53 -3262
rect -1 -3422 139 -3262
rect 191 -3422 331 -3262
rect 383 -3422 523 -3262
rect 844 -3422 907 -3262
rect 959 -3422 1099 -3262
rect 1151 -3422 1164 -3262
rect -1226 -3640 524 -3422
rect 844 -3640 1164 -3422
rect -1226 -3800 -1205 -3640
rect -1153 -3800 -1013 -3640
rect -961 -3800 -821 -3640
rect -769 -3800 -629 -3640
rect -577 -3800 -437 -3640
rect -385 -3800 -245 -3640
rect -193 -3800 -53 -3640
rect -1 -3800 139 -3640
rect 191 -3800 331 -3640
rect 383 -3800 523 -3640
rect 844 -3800 907 -3640
rect 959 -3800 1099 -3640
rect 1151 -3800 1164 -3640
rect -1205 -3810 -1153 -3800
rect -1013 -3810 -961 -3800
rect -821 -3810 -769 -3800
rect -629 -3810 -577 -3800
rect -437 -3810 -385 -3800
rect -245 -3810 -193 -3800
rect -53 -3810 -1 -3800
rect 139 -3810 191 -3800
rect 331 -3810 383 -3800
rect 523 -3810 844 -3800
rect 907 -3810 959 -3800
rect 1099 -3810 1151 -3800
rect -146 -3870 174 -3860
rect 1244 -3870 1384 -3192
rect -1116 -3880 -146 -3870
rect 174 -3880 1384 -3870
rect -1380 -4020 -1270 -4010
rect -1116 -4040 -1109 -3880
rect -1057 -4040 -917 -3880
rect -865 -4040 -725 -3880
rect -673 -4040 -533 -3880
rect -481 -4040 -341 -3880
rect -289 -4040 -149 -3880
rect 174 -4040 235 -3880
rect 287 -4040 427 -3880
rect 479 -4040 619 -3880
rect 671 -4040 811 -3880
rect 863 -4040 1003 -3880
rect 1055 -4040 1195 -3880
rect 1247 -4040 1384 -3880
rect -1116 -4050 -146 -4040
rect 174 -4050 1384 -4040
rect -146 -4060 174 -4050
rect -1380 -8760 -1270 -4120
rect -1087 -4520 -1035 -4515
rect -891 -4520 -839 -4515
rect -695 -4520 -643 -4515
rect -499 -4520 -447 -4515
rect -303 -4520 -251 -4515
rect -107 -4520 -55 -4515
rect 89 -4520 141 -4515
rect 285 -4520 337 -4515
rect 711 -4520 763 -4515
rect 907 -4520 959 -4515
rect 1103 -4520 1155 -4515
rect 1299 -4520 1351 -4515
rect 1495 -4520 1547 -4515
rect 1691 -4520 1743 -4515
rect 1887 -4520 1939 -4515
rect 2083 -4520 2135 -4515
rect -1096 -4525 2304 -4520
rect -1096 -4685 -1087 -4525
rect -1035 -4685 -891 -4525
rect -839 -4685 -695 -4525
rect -643 -4685 -499 -4525
rect -447 -4685 -303 -4525
rect -251 -4685 -107 -4525
rect -55 -4685 89 -4525
rect 141 -4685 285 -4525
rect 337 -4540 711 -4525
rect 337 -4680 354 -4540
rect 594 -4680 711 -4540
rect 337 -4685 711 -4680
rect 763 -4685 907 -4525
rect 959 -4685 1103 -4525
rect 1155 -4685 1299 -4525
rect 1351 -4685 1495 -4525
rect 1547 -4685 1691 -4525
rect 1743 -4685 1887 -4525
rect 1939 -4685 2083 -4525
rect 2135 -4685 2304 -4525
rect -1096 -4690 2304 -4685
rect -1087 -4695 -1035 -4690
rect -891 -4695 -839 -4690
rect -695 -4695 -643 -4690
rect -499 -4695 -447 -4690
rect -303 -4695 -251 -4690
rect -107 -4695 -55 -4690
rect 89 -4695 141 -4690
rect 285 -4695 337 -4690
rect 711 -4695 763 -4690
rect 907 -4695 959 -4690
rect 1103 -4695 1155 -4690
rect 1299 -4695 1351 -4690
rect 1495 -4695 1547 -4690
rect 1691 -4695 1743 -4690
rect 1887 -4695 1939 -4690
rect 2054 -4700 2304 -4690
rect -1185 -4760 -1133 -4755
rect -989 -4760 -937 -4755
rect -793 -4760 -741 -4755
rect -597 -4760 -545 -4755
rect -401 -4760 -349 -4755
rect -205 -4760 -153 -4755
rect -9 -4760 43 -4755
rect 187 -4760 239 -4755
rect 613 -4760 665 -4755
rect 809 -4760 861 -4755
rect 1005 -4760 1057 -4755
rect 1201 -4760 1253 -4755
rect 1397 -4760 1449 -4755
rect 1593 -4760 1645 -4755
rect 1789 -4760 1841 -4755
rect 1985 -4760 2037 -4755
rect -1196 -4765 2044 -4760
rect -1196 -4925 -1185 -4765
rect -1133 -4925 -989 -4765
rect -937 -4925 -793 -4765
rect -741 -4925 -597 -4765
rect -545 -4925 -401 -4765
rect -349 -4925 -205 -4765
rect -153 -4925 -9 -4765
rect 43 -4925 187 -4765
rect 239 -4925 613 -4765
rect 665 -4925 809 -4765
rect 861 -4770 1005 -4765
rect 1057 -4770 1201 -4765
rect 1253 -4770 1397 -4765
rect 861 -4920 974 -4770
rect 1374 -4920 1397 -4770
rect 861 -4925 1005 -4920
rect 1057 -4925 1201 -4920
rect 1253 -4925 1397 -4920
rect 1449 -4925 1593 -4765
rect 1645 -4925 1789 -4765
rect 1841 -4925 1985 -4765
rect 2037 -4925 2044 -4765
rect -1196 -4930 2044 -4925
rect -1185 -4935 -1133 -4930
rect -989 -4935 -937 -4930
rect -793 -4935 -741 -4930
rect -597 -4935 -545 -4930
rect -401 -4935 -349 -4930
rect -205 -4935 -153 -4930
rect -9 -4935 43 -4930
rect 187 -4935 239 -4930
rect 613 -4935 665 -4930
rect 809 -4935 861 -4930
rect 1005 -4935 1057 -4930
rect 1201 -4935 1253 -4930
rect 1397 -4935 1449 -4930
rect 1593 -4935 1645 -4930
rect 1789 -4935 1841 -4930
rect 1985 -4935 2037 -4930
rect 2164 -4980 2304 -4700
rect 2164 -5000 3894 -4980
rect -1185 -5160 -1133 -5151
rect -989 -5160 -937 -5151
rect -793 -5160 -741 -5151
rect -597 -5160 -545 -5151
rect -401 -5160 -349 -5151
rect -205 -5160 -153 -5151
rect -9 -5160 43 -5151
rect 187 -5160 239 -5151
rect 613 -5160 665 -5151
rect 809 -5160 861 -5151
rect 1005 -5160 1057 -5151
rect 1201 -5160 1253 -5151
rect 1397 -5160 1449 -5151
rect 1593 -5160 1645 -5151
rect 1789 -5160 1841 -5151
rect 1985 -5160 2037 -5151
rect -1196 -5161 2044 -5160
rect -1196 -5321 -1185 -5161
rect -1133 -5321 -989 -5161
rect -937 -5321 -793 -5161
rect -741 -5321 -597 -5161
rect -545 -5321 -401 -5161
rect -349 -5321 -205 -5161
rect -153 -5321 -9 -5161
rect 43 -5321 187 -5161
rect 239 -5321 613 -5161
rect 665 -5321 809 -5161
rect 861 -5170 1005 -5161
rect 1057 -5170 1201 -5161
rect 1253 -5170 1397 -5161
rect 861 -5320 984 -5170
rect 1384 -5320 1397 -5170
rect 861 -5321 1005 -5320
rect 1057 -5321 1201 -5320
rect 1253 -5321 1397 -5320
rect 1449 -5321 1593 -5161
rect 1645 -5321 1789 -5161
rect 1841 -5321 1985 -5161
rect 2037 -5321 2044 -5161
rect -1196 -5330 2044 -5321
rect -1185 -5331 -1133 -5330
rect -989 -5331 -937 -5330
rect -793 -5331 -741 -5330
rect -597 -5331 -545 -5330
rect -401 -5331 -349 -5330
rect -205 -5331 -153 -5330
rect -9 -5331 43 -5330
rect 187 -5331 239 -5330
rect 613 -5331 665 -5330
rect 809 -5331 861 -5330
rect 1005 -5331 1057 -5330
rect 1201 -5331 1253 -5330
rect 1397 -5331 1449 -5330
rect 1593 -5331 1645 -5330
rect 1789 -5331 1841 -5330
rect 1985 -5331 2037 -5330
rect 2164 -5390 2214 -5000
rect -1087 -5400 -1035 -5391
rect -891 -5400 -839 -5391
rect -695 -5400 -643 -5391
rect -499 -5400 -447 -5391
rect -303 -5400 -251 -5391
rect -107 -5400 -55 -5391
rect 89 -5400 141 -5391
rect 285 -5400 337 -5391
rect 711 -5400 763 -5391
rect 907 -5400 959 -5391
rect 1103 -5400 1155 -5391
rect 1299 -5400 1351 -5391
rect 1495 -5400 1547 -5391
rect 1691 -5400 1743 -5391
rect 1887 -5400 1939 -5391
rect 2054 -5400 2214 -5390
rect -1087 -5401 2214 -5400
rect -1035 -5560 -891 -5401
rect -1087 -5571 -1035 -5561
rect -839 -5560 -695 -5401
rect -891 -5571 -839 -5561
rect -643 -5560 -499 -5401
rect -695 -5571 -643 -5561
rect -447 -5560 -303 -5401
rect -499 -5571 -447 -5561
rect -251 -5560 -107 -5401
rect -303 -5571 -251 -5561
rect -55 -5560 89 -5401
rect -107 -5571 -55 -5561
rect 141 -5560 285 -5401
rect 89 -5571 141 -5561
rect 337 -5420 711 -5401
rect 337 -5560 354 -5420
rect 594 -5560 711 -5420
rect 337 -5561 614 -5560
rect 285 -5571 614 -5561
rect 763 -5560 907 -5401
rect 711 -5571 763 -5561
rect 959 -5560 1103 -5401
rect 907 -5571 959 -5561
rect 1155 -5560 1299 -5401
rect 1103 -5571 1155 -5561
rect 1351 -5560 1495 -5401
rect 1299 -5571 1351 -5561
rect 1547 -5560 1691 -5401
rect 1495 -5571 1547 -5561
rect 1743 -5560 1887 -5401
rect 1691 -5571 1743 -5561
rect 1939 -5560 2083 -5401
rect 1887 -5571 1939 -5561
rect 2135 -5560 2214 -5401
rect 2344 -5177 3894 -5000
rect 2344 -5337 2573 -5177
rect 2625 -5337 2889 -5177
rect 2941 -5337 3205 -5177
rect 3257 -5337 3521 -5177
rect 3573 -5337 3837 -5177
rect 3889 -5260 3894 -5177
rect 4190 -5080 4290 -5070
rect 5080 -5080 5170 -5070
rect 4290 -5200 5080 -5080
rect 4190 -5210 4290 -5200
rect 5080 -5210 5170 -5200
rect 3889 -5337 4500 -5260
rect 2344 -5340 4500 -5337
rect 2573 -5347 2625 -5340
rect 2889 -5347 2941 -5340
rect 3205 -5347 3257 -5340
rect 3521 -5347 3573 -5340
rect 3837 -5347 3889 -5340
rect 2834 -5400 3274 -5390
rect 2415 -5410 2467 -5407
rect 2731 -5410 2783 -5407
rect 2083 -5571 2135 -5561
rect 2214 -5570 2344 -5560
rect 2414 -5417 2834 -5410
rect 3363 -5410 3415 -5407
rect 3679 -5410 3731 -5407
rect 3995 -5410 4047 -5407
rect 3274 -5417 4054 -5410
rect 314 -5580 614 -5571
rect 2414 -5577 2415 -5417
rect 2467 -5577 2731 -5417
rect 2783 -5577 2834 -5417
rect 3274 -5577 3363 -5417
rect 3415 -5577 3679 -5417
rect 3731 -5577 3995 -5417
rect 4047 -5577 4054 -5417
rect 2414 -5580 2834 -5577
rect 3274 -5580 4054 -5577
rect 2415 -5587 2467 -5580
rect 2731 -5587 2783 -5580
rect 2834 -5590 3274 -5580
rect 3363 -5587 3415 -5580
rect 3679 -5587 3731 -5580
rect 3995 -5587 4047 -5580
rect 524 -5982 844 -5980
rect -1087 -5990 -1035 -5982
rect -891 -5990 -839 -5982
rect -695 -5990 -643 -5982
rect -499 -5990 -447 -5982
rect -303 -5990 -251 -5982
rect -107 -5990 -55 -5982
rect 89 -5990 141 -5982
rect 285 -5990 337 -5982
rect 481 -5990 844 -5982
rect 873 -5990 925 -5982
rect 1069 -5990 1121 -5982
rect 1265 -5990 1317 -5982
rect -1096 -5992 524 -5990
rect 844 -5992 1324 -5990
rect -1096 -6152 -1087 -5992
rect -1035 -6152 -891 -5992
rect -839 -6152 -695 -5992
rect -643 -6152 -499 -5992
rect -447 -6152 -303 -5992
rect -251 -6152 -107 -5992
rect -55 -6152 89 -5992
rect 141 -6152 285 -5992
rect 337 -6152 481 -5992
rect 844 -6152 873 -5992
rect 925 -6152 1069 -5992
rect 1121 -6152 1265 -5992
rect 1317 -6152 1324 -5992
rect -1096 -6160 524 -6152
rect 844 -6160 1324 -6152
rect -1087 -6162 -1035 -6160
rect -891 -6162 -839 -6160
rect -695 -6162 -643 -6160
rect -499 -6162 -447 -6160
rect -303 -6162 -251 -6160
rect -107 -6162 -55 -6160
rect 89 -6162 141 -6160
rect 285 -6162 337 -6160
rect 481 -6162 844 -6160
rect 873 -6162 925 -6160
rect 1069 -6162 1121 -6160
rect 1265 -6162 1317 -6160
rect 524 -6170 844 -6162
rect 2164 -6220 2414 -6210
rect -1185 -6230 -1133 -6222
rect -989 -6230 -937 -6222
rect -793 -6230 -741 -6222
rect -597 -6230 -545 -6222
rect -401 -6230 -349 -6222
rect -205 -6230 -153 -6222
rect -9 -6230 43 -6222
rect 187 -6230 239 -6222
rect 383 -6230 435 -6222
rect 579 -6230 631 -6222
rect 775 -6230 827 -6222
rect 971 -6230 1023 -6222
rect 1167 -6230 1219 -6222
rect -1186 -6232 2164 -6230
rect -1186 -6392 -1185 -6232
rect -1133 -6392 -989 -6232
rect -937 -6392 -793 -6232
rect -741 -6392 -597 -6232
rect -545 -6392 -401 -6232
rect -349 -6392 -205 -6232
rect -153 -6392 -9 -6232
rect 43 -6392 187 -6232
rect 239 -6392 383 -6232
rect 435 -6392 579 -6232
rect 631 -6392 775 -6232
rect 827 -6392 971 -6232
rect 1023 -6240 1167 -6232
rect 1219 -6240 2164 -6232
rect 1384 -6390 2164 -6240
rect 1023 -6392 1167 -6390
rect 1219 -6392 2164 -6390
rect -1186 -6400 2164 -6392
rect -1185 -6402 -1133 -6400
rect -989 -6402 -937 -6400
rect -793 -6402 -741 -6400
rect -597 -6402 -545 -6400
rect -401 -6402 -349 -6400
rect -205 -6402 -153 -6400
rect -9 -6402 43 -6400
rect 187 -6402 239 -6400
rect 383 -6402 435 -6400
rect 579 -6402 631 -6400
rect 775 -6402 827 -6400
rect 971 -6402 1023 -6400
rect 1167 -6402 1219 -6400
rect 2834 -6300 3274 -6290
rect 2164 -6420 2414 -6410
rect 2464 -6312 2834 -6300
rect 3274 -6312 3914 -6300
rect 2464 -6472 2475 -6312
rect 2527 -6472 2671 -6312
rect 2723 -6472 2834 -6312
rect 3311 -6472 3455 -6312
rect 3507 -6472 3651 -6312
rect 3703 -6472 3847 -6312
rect 3899 -6472 3914 -6312
rect 2464 -6480 2834 -6472
rect 3274 -6480 3914 -6472
rect 2475 -6482 2527 -6480
rect 2671 -6482 2723 -6480
rect 2834 -6482 3311 -6480
rect 3455 -6482 3507 -6480
rect 3651 -6482 3703 -6480
rect 3847 -6482 3899 -6480
rect 2834 -6490 3274 -6482
rect 2564 -6552 4114 -6540
rect -1186 -6610 1384 -6600
rect -1186 -6770 -1185 -6610
rect -1133 -6770 -989 -6610
rect -937 -6770 -793 -6610
rect -741 -6770 -597 -6610
rect -545 -6770 -401 -6610
rect -349 -6770 -205 -6610
rect -153 -6770 -9 -6610
rect 43 -6770 187 -6610
rect 239 -6770 383 -6610
rect 435 -6770 579 -6610
rect 631 -6770 775 -6610
rect 827 -6770 971 -6610
rect 2564 -6712 2573 -6552
rect 2625 -6712 2769 -6552
rect 2821 -6712 2965 -6552
rect 3017 -6712 3161 -6552
rect 3213 -6712 3357 -6552
rect 3409 -6712 3553 -6552
rect 3605 -6712 3749 -6552
rect 3801 -6712 3945 -6552
rect 3997 -6712 4114 -6552
rect 2564 -6720 4114 -6712
rect 2573 -6722 2734 -6720
rect 2769 -6722 2821 -6720
rect 2965 -6722 3017 -6720
rect 3161 -6722 3213 -6720
rect 3357 -6722 3409 -6720
rect 3553 -6722 3605 -6720
rect 3749 -6722 3801 -6720
rect 1023 -6770 1167 -6760
rect 1219 -6770 1384 -6760
rect 1454 -6750 1684 -6740
rect 2204 -6750 2284 -6740
rect 2574 -6750 2734 -6722
rect 3924 -6730 4174 -6720
rect -1185 -6780 -1133 -6770
rect -989 -6780 -937 -6770
rect -793 -6780 -741 -6770
rect -597 -6780 -545 -6770
rect -401 -6780 -349 -6770
rect -205 -6780 -153 -6770
rect -9 -6780 43 -6770
rect 187 -6780 239 -6770
rect 383 -6780 435 -6770
rect 579 -6780 631 -6770
rect 775 -6780 827 -6770
rect 971 -6780 1023 -6770
rect 1167 -6780 1219 -6770
rect -1087 -6850 -1035 -6840
rect -891 -6850 -839 -6840
rect -695 -6850 -643 -6840
rect -499 -6850 -447 -6840
rect -303 -6850 -251 -6840
rect -107 -6850 -55 -6840
rect 89 -6850 141 -6840
rect 285 -6850 337 -6840
rect 424 -6850 1317 -6840
rect -1096 -7010 -1087 -6850
rect -1035 -7010 -891 -6850
rect -839 -7010 -695 -6850
rect -643 -7010 -499 -6850
rect -447 -7010 -303 -6850
rect -251 -7010 -107 -6850
rect -55 -7010 89 -6850
rect 141 -7010 285 -6850
rect 337 -7010 481 -6850
rect 844 -7010 873 -6850
rect 925 -7010 1069 -6850
rect 1121 -7010 1265 -6850
rect 1317 -7010 1324 -6850
rect 1684 -6910 2204 -6750
rect 2284 -6910 2734 -6750
rect 1454 -6920 1684 -6910
rect 2204 -6920 2284 -6910
rect 2564 -6920 2734 -6910
rect 4004 -6920 4054 -6730
rect -1096 -7436 524 -7010
rect 844 -7436 1324 -7010
rect 2564 -6930 4054 -6920
rect 2564 -7090 2573 -6930
rect 2625 -7090 2769 -6930
rect 2821 -7090 2965 -6930
rect 3017 -7090 3161 -6930
rect 3213 -7090 3357 -6930
rect 3409 -7090 3553 -6930
rect 3605 -7090 3749 -6930
rect 3801 -7090 3945 -6930
rect 3997 -6940 4054 -6930
rect 3997 -6950 4174 -6940
rect 3997 -7090 4114 -6950
rect 2564 -7100 4114 -7090
rect 2834 -7160 3274 -7150
rect 2464 -7170 2834 -7160
rect 3274 -7170 3914 -7160
rect 2464 -7330 2475 -7170
rect 2527 -7330 2671 -7170
rect 2723 -7330 2834 -7170
rect 3311 -7330 3455 -7170
rect 3507 -7330 3651 -7170
rect 3703 -7330 3847 -7170
rect 3899 -7330 3914 -7170
rect 2464 -7340 2834 -7330
rect 3274 -7340 3914 -7330
rect 2834 -7350 3274 -7340
rect -1096 -7596 -1087 -7436
rect -1035 -7596 -891 -7436
rect -839 -7596 -695 -7436
rect -643 -7596 -499 -7436
rect -447 -7596 -303 -7436
rect -251 -7596 -107 -7436
rect -55 -7596 89 -7436
rect 141 -7596 285 -7436
rect 337 -7596 481 -7436
rect 844 -7596 873 -7436
rect 925 -7596 1069 -7436
rect 1121 -7596 1265 -7436
rect 1317 -7596 1324 -7436
rect -1096 -7600 524 -7596
rect 844 -7600 1324 -7596
rect 4320 -7540 4500 -5340
rect -1087 -7606 -1035 -7600
rect -891 -7606 -839 -7600
rect -695 -7606 -643 -7600
rect -499 -7606 -447 -7600
rect -303 -7606 -251 -7600
rect -107 -7606 -55 -7600
rect 89 -7606 141 -7600
rect 285 -7606 337 -7600
rect 434 -7606 925 -7600
rect 1069 -7606 1121 -7600
rect 1265 -7606 1317 -7600
rect 434 -7610 924 -7606
rect -1185 -7670 -1133 -7666
rect -989 -7670 -937 -7666
rect -793 -7670 -741 -7666
rect -597 -7670 -545 -7666
rect -401 -7670 -349 -7666
rect -205 -7670 -153 -7666
rect -9 -7670 43 -7666
rect 187 -7670 239 -7666
rect 383 -7670 435 -7666
rect 579 -7670 631 -7666
rect 775 -7670 827 -7666
rect 971 -7670 1023 -7666
rect 1167 -7670 1219 -7666
rect -1196 -7676 1384 -7670
rect -1196 -7836 -1185 -7676
rect -1133 -7836 -989 -7676
rect -937 -7836 -793 -7676
rect -741 -7836 -597 -7676
rect -545 -7836 -401 -7676
rect -349 -7836 -205 -7676
rect -153 -7836 -9 -7676
rect 43 -7836 187 -7676
rect 239 -7836 383 -7676
rect 435 -7836 579 -7676
rect 631 -7836 775 -7676
rect 827 -7836 971 -7676
rect 1023 -7680 1167 -7676
rect 1219 -7680 1384 -7676
rect 4320 -7710 5050 -7540
rect 1023 -7836 1167 -7830
rect 1219 -7836 1384 -7830
rect -1196 -7840 1384 -7836
rect -1185 -7846 -1133 -7840
rect -989 -7846 -937 -7840
rect -793 -7846 -741 -7840
rect -597 -7846 -545 -7840
rect -401 -7846 -349 -7840
rect -205 -7846 -153 -7840
rect -9 -7846 43 -7840
rect 187 -7846 239 -7840
rect 383 -7846 435 -7840
rect 579 -7846 631 -7840
rect 775 -7846 827 -7840
rect 971 -7846 1023 -7840
rect 1167 -7846 1219 -7840
rect 2850 -7990 3020 -7980
rect -1186 -8050 1804 -8040
rect -1186 -8054 984 -8050
rect -1186 -8210 -1185 -8054
rect -1133 -8210 -989 -8054
rect -1185 -8224 -1133 -8214
rect -937 -8210 -793 -8054
rect -989 -8224 -937 -8214
rect -741 -8210 -597 -8054
rect -793 -8224 -741 -8214
rect -545 -8210 -401 -8054
rect -597 -8224 -545 -8214
rect -349 -8210 -205 -8054
rect -401 -8224 -349 -8214
rect -153 -8210 -9 -8054
rect -205 -8224 -153 -8214
rect 43 -8210 187 -8054
rect -9 -8224 43 -8214
rect 239 -8210 383 -8054
rect 187 -8224 239 -8214
rect 435 -8210 579 -8054
rect 383 -8224 435 -8214
rect 631 -8210 775 -8054
rect 579 -8224 631 -8214
rect 827 -8210 971 -8054
rect 1384 -8080 1804 -8050
rect 1384 -8090 2724 -8080
rect 1384 -8200 1701 -8090
rect 775 -8224 827 -8214
rect 1023 -8210 1167 -8200
rect 971 -8224 1023 -8214
rect 1219 -8210 1701 -8200
rect 1167 -8224 1219 -8214
rect 1694 -8250 1701 -8210
rect 1753 -8250 1893 -8090
rect 1945 -8250 2085 -8090
rect 2137 -8250 2277 -8090
rect 2329 -8250 2469 -8090
rect 2521 -8250 2661 -8090
rect 2713 -8250 2724 -8090
rect 2850 -8150 3020 -8140
rect 3590 -8090 4620 -8080
rect 1694 -8260 2724 -8250
rect 3590 -8250 3597 -8090
rect 3649 -8250 3789 -8090
rect 3841 -8250 3981 -8090
rect 4033 -8250 4173 -8090
rect 4225 -8250 4365 -8090
rect 4417 -8250 4550 -8090
rect 3590 -8260 4620 -8250
rect 524 -8284 844 -8280
rect -1087 -8290 -1035 -8284
rect -891 -8290 -839 -8284
rect -695 -8290 -643 -8284
rect -499 -8290 -447 -8284
rect -303 -8290 -251 -8284
rect -107 -8290 -55 -8284
rect 89 -8290 141 -8284
rect 285 -8290 337 -8284
rect 481 -8290 844 -8284
rect 873 -8290 925 -8284
rect 1069 -8290 1121 -8284
rect 1265 -8290 1317 -8284
rect -1096 -8294 524 -8290
rect 844 -8294 1324 -8290
rect -1096 -8454 -1087 -8294
rect -1035 -8454 -891 -8294
rect -839 -8454 -695 -8294
rect -643 -8454 -499 -8294
rect -447 -8454 -303 -8294
rect -251 -8454 -107 -8294
rect -55 -8454 89 -8294
rect 141 -8454 285 -8294
rect 337 -8454 481 -8294
rect 844 -8454 873 -8294
rect 925 -8454 1069 -8294
rect 1121 -8454 1265 -8294
rect 1317 -8454 1324 -8294
rect -1096 -8460 524 -8454
rect 844 -8460 1324 -8454
rect 1604 -8330 2954 -8320
rect -1087 -8464 -1035 -8460
rect -891 -8464 -839 -8460
rect -695 -8464 -643 -8460
rect -499 -8464 -447 -8460
rect -303 -8464 -251 -8460
rect -107 -8464 -55 -8460
rect 89 -8464 141 -8460
rect 285 -8464 337 -8460
rect 481 -8464 844 -8460
rect 873 -8464 925 -8460
rect 1069 -8464 1121 -8460
rect 1265 -8464 1317 -8460
rect 524 -8470 844 -8464
rect 1604 -8490 1605 -8330
rect 1657 -8490 1797 -8330
rect 1849 -8490 1989 -8330
rect 2041 -8490 2181 -8330
rect 2233 -8490 2373 -8330
rect 2425 -8490 2565 -8330
rect 2617 -8490 2757 -8330
rect 2809 -8490 2954 -8330
rect 1604 -8500 2954 -8490
rect 3500 -8330 4850 -8320
rect 3500 -8490 3501 -8330
rect 3553 -8490 3693 -8330
rect 3745 -8490 3885 -8330
rect 3937 -8490 4077 -8330
rect 4129 -8490 4269 -8330
rect 4321 -8490 4461 -8330
rect 4513 -8490 4653 -8330
rect 4705 -8490 4850 -8330
rect 3500 -8500 4850 -8490
rect -146 -8840 174 -8830
rect -1109 -8850 -1057 -8846
rect -917 -8850 -865 -8846
rect -725 -8850 -673 -8846
rect -533 -8850 -481 -8846
rect -341 -8850 -289 -8846
rect -149 -8850 -146 -8846
rect -1380 -8860 -1270 -8850
rect -1116 -8856 -146 -8850
rect 235 -8850 287 -8846
rect 427 -8850 479 -8846
rect 619 -8850 671 -8846
rect 811 -8850 863 -8846
rect 1003 -8850 1055 -8846
rect 1195 -8850 1247 -8846
rect 174 -8856 1384 -8850
rect -1116 -9016 -1109 -8856
rect -1057 -9016 -917 -8856
rect -865 -9016 -725 -8856
rect -673 -9016 -533 -8856
rect -481 -9016 -341 -8856
rect -289 -9016 -149 -8856
rect 174 -9016 235 -8856
rect 287 -9016 427 -8856
rect 479 -9016 619 -8856
rect 671 -9016 811 -8856
rect 863 -9016 1003 -8856
rect 1055 -9016 1195 -8856
rect 1247 -9016 1384 -8856
rect 2654 -8880 2954 -8500
rect 4550 -8880 4850 -8500
rect 4930 -8540 5050 -7710
rect 4930 -8650 6350 -8540
rect -1116 -9020 -146 -9016
rect 174 -9020 1384 -9016
rect -1109 -9026 -1057 -9020
rect -917 -9026 -865 -9020
rect -725 -9026 -673 -9020
rect -533 -9026 -481 -9020
rect -341 -9026 -289 -9020
rect -149 -9026 174 -9020
rect 235 -9026 287 -9020
rect 427 -9026 479 -9020
rect 619 -9026 671 -9020
rect 811 -9026 863 -9020
rect 1003 -9026 1055 -9020
rect 1195 -9026 1384 -9020
rect -146 -9030 174 -9026
rect -1205 -9090 -1153 -9086
rect -1013 -9090 -961 -9086
rect -821 -9090 -769 -9086
rect -629 -9090 -577 -9086
rect -437 -9090 -385 -9086
rect -245 -9090 -193 -9086
rect -53 -9090 -1 -9086
rect 139 -9090 191 -9086
rect 331 -9090 383 -9086
rect 523 -9090 575 -9086
rect 715 -9090 767 -9086
rect 907 -9090 959 -9086
rect 1099 -9090 1151 -9086
rect -1216 -9096 1154 -9090
rect -1216 -9256 -1205 -9096
rect -1153 -9256 -1013 -9096
rect -961 -9256 -821 -9096
rect -769 -9256 -629 -9096
rect -577 -9256 -437 -9096
rect -385 -9256 -245 -9096
rect -193 -9256 -53 -9096
rect -1 -9256 139 -9096
rect 191 -9256 331 -9096
rect 383 -9256 523 -9096
rect 575 -9100 715 -9096
rect 767 -9100 907 -9096
rect 844 -9256 907 -9100
rect 959 -9256 1099 -9096
rect 1151 -9256 1154 -9096
rect -1216 -9474 524 -9256
rect 844 -9474 1154 -9256
rect -1216 -9634 -1205 -9474
rect -1153 -9634 -1013 -9474
rect -961 -9634 -821 -9474
rect -769 -9634 -629 -9474
rect -577 -9634 -437 -9474
rect -385 -9634 -245 -9474
rect -193 -9634 -53 -9474
rect -1 -9634 139 -9474
rect 191 -9634 331 -9474
rect 383 -9634 523 -9474
rect 844 -9634 907 -9474
rect 959 -9634 1099 -9474
rect 1151 -9634 1154 -9474
rect -1216 -9640 524 -9634
rect 844 -9640 1154 -9634
rect 1244 -9130 1384 -9026
rect 1844 -8910 2954 -8880
rect 1844 -9070 1863 -8910
rect 1915 -9070 2379 -8910
rect 2431 -9070 2895 -8910
rect 2947 -9070 2954 -8910
rect 1844 -9080 2954 -9070
rect 3740 -8910 4850 -8880
rect 3740 -9070 3759 -8910
rect 3811 -9070 4275 -8910
rect 4327 -9070 4791 -8910
rect 4843 -9070 4850 -8910
rect 3740 -9080 4850 -9070
rect 5440 -8910 5500 -8900
rect 5640 -8910 5700 -8900
rect 5830 -8910 5890 -8900
rect 5500 -9090 5640 -8910
rect 5700 -9090 5830 -8910
rect 5440 -9100 5500 -9090
rect 5640 -9100 5700 -9090
rect 5830 -9100 5890 -9090
rect 1244 -9140 1474 -9130
rect 1244 -9210 1344 -9140
rect 1474 -9150 5110 -9140
rect 5540 -9150 5600 -9140
rect 5740 -9150 5800 -9140
rect 5930 -9150 5990 -9140
rect 1474 -9210 1605 -9150
rect -1205 -9644 -1153 -9640
rect -1013 -9644 -961 -9640
rect -821 -9644 -769 -9640
rect -629 -9644 -577 -9640
rect -437 -9644 -385 -9640
rect -245 -9644 -193 -9640
rect -53 -9644 -1 -9640
rect 139 -9644 191 -9640
rect 331 -9644 383 -9640
rect 523 -9644 844 -9640
rect 907 -9644 959 -9640
rect 1099 -9644 1151 -9640
rect 524 -9650 844 -9644
rect 1244 -9650 1250 -9210
rect 1480 -9310 1605 -9210
rect 1657 -9310 2121 -9150
rect 2173 -9310 2637 -9150
rect 2689 -9310 3153 -9150
rect 3205 -9310 3501 -9150
rect 3553 -9310 4017 -9150
rect 4069 -9310 4533 -9150
rect 4585 -9310 5049 -9150
rect 5101 -9310 5540 -9150
rect 5600 -9310 5740 -9150
rect 5800 -9310 5930 -9150
rect 1480 -9320 3214 -9310
rect 3490 -9320 5110 -9310
rect 5540 -9320 5600 -9310
rect 5740 -9320 5800 -9310
rect 5930 -9320 5990 -9310
rect 6060 -9300 6130 -9290
rect 6060 -9420 6130 -9410
rect 1244 -9660 1480 -9650
rect 1244 -9704 1384 -9660
rect -1109 -9710 -1057 -9704
rect -917 -9710 -865 -9704
rect -725 -9710 -673 -9704
rect -533 -9710 -481 -9704
rect -341 -9710 -289 -9704
rect -149 -9710 -97 -9704
rect 43 -9710 95 -9704
rect 235 -9710 287 -9704
rect 427 -9710 479 -9704
rect 619 -9710 671 -9704
rect 811 -9710 863 -9704
rect 1003 -9710 1055 -9704
rect 1195 -9710 1384 -9704
rect -1116 -9714 1384 -9710
rect -1116 -9874 -1109 -9714
rect -1057 -9874 -917 -9714
rect -865 -9874 -725 -9714
rect -673 -9874 -533 -9714
rect -481 -9874 -341 -9714
rect -289 -9874 -149 -9714
rect -97 -9720 43 -9714
rect 95 -9720 235 -9714
rect 174 -9874 235 -9720
rect 287 -9874 427 -9714
rect 479 -9874 619 -9714
rect 671 -9874 811 -9714
rect 863 -9874 1003 -9714
rect 1055 -9874 1195 -9714
rect 1247 -9874 1384 -9714
rect 6230 -9700 6350 -8650
rect 6230 -9810 6760 -9700
rect -1116 -10092 -146 -9874
rect 174 -10092 1384 -9874
rect 6390 -9960 6460 -9950
rect 6390 -10080 6460 -10070
rect -1116 -10252 -1109 -10092
rect -1057 -10252 -917 -10092
rect -865 -10252 -725 -10092
rect -673 -10252 -533 -10092
rect -481 -10252 -341 -10092
rect -289 -10252 -149 -10092
rect 174 -10252 235 -10092
rect 287 -10252 427 -10092
rect 479 -10252 619 -10092
rect 671 -10252 811 -10092
rect 863 -10252 1003 -10092
rect 1055 -10252 1195 -10092
rect 1247 -10252 1384 -10092
rect -1116 -10260 -146 -10252
rect 174 -10260 1384 -10252
rect -1109 -10262 -1057 -10260
rect -917 -10262 -865 -10260
rect -725 -10262 -673 -10260
rect -533 -10262 -481 -10260
rect -341 -10262 -289 -10260
rect -149 -10262 174 -10260
rect 235 -10262 287 -10260
rect 427 -10262 479 -10260
rect 619 -10262 671 -10260
rect 811 -10262 863 -10260
rect 1003 -10262 1055 -10260
rect 1195 -10262 1384 -10260
rect -146 -10270 174 -10262
rect -1226 -10330 1164 -10320
rect -1226 -10332 524 -10330
rect 844 -10332 1164 -10330
rect -1226 -10492 -1205 -10332
rect -1153 -10492 -1013 -10332
rect -961 -10492 -821 -10332
rect -769 -10492 -629 -10332
rect -577 -10492 -437 -10332
rect -385 -10492 -245 -10332
rect -193 -10492 -53 -10332
rect -1 -10492 139 -10332
rect 191 -10492 331 -10332
rect 383 -10492 523 -10332
rect 844 -10492 907 -10332
rect 959 -10492 1099 -10332
rect 1151 -10492 1164 -10332
rect -1226 -10710 524 -10492
rect 844 -10710 1164 -10492
rect -1226 -10870 -1205 -10710
rect -1153 -10870 -1013 -10710
rect -961 -10870 -821 -10710
rect -769 -10870 -629 -10710
rect -577 -10870 -437 -10710
rect -385 -10870 -245 -10710
rect -193 -10870 -53 -10710
rect -1 -10870 139 -10710
rect 191 -10870 331 -10710
rect 383 -10870 523 -10710
rect 844 -10870 907 -10710
rect 959 -10870 1099 -10710
rect 1151 -10870 1164 -10710
rect -1205 -10880 -1153 -10870
rect -1013 -10880 -961 -10870
rect -821 -10880 -769 -10870
rect -629 -10880 -577 -10870
rect -437 -10880 -385 -10870
rect -245 -10880 -193 -10870
rect -53 -10880 -1 -10870
rect 139 -10880 191 -10870
rect 331 -10880 383 -10870
rect 523 -10880 844 -10870
rect 907 -10880 959 -10870
rect 1099 -10880 1151 -10870
rect -146 -10940 174 -10930
rect 1244 -10940 1384 -10262
rect 6620 -10200 6760 -9810
rect 6620 -10330 6760 -10320
rect -1116 -10950 -146 -10940
rect 174 -10950 1384 -10940
rect -1116 -11110 -1109 -10950
rect -1057 -11110 -917 -10950
rect -865 -11110 -725 -10950
rect -673 -11110 -533 -10950
rect -481 -11110 -341 -10950
rect -289 -11110 -149 -10950
rect 174 -11110 235 -10950
rect 287 -11110 427 -10950
rect 479 -11110 619 -10950
rect 671 -11110 811 -10950
rect 863 -11110 1003 -10950
rect 1055 -11110 1195 -10950
rect 1247 -11110 1384 -10950
rect -1116 -11120 -146 -11110
rect 174 -11120 1384 -11110
rect -146 -11130 174 -11120
<< via2 >>
rect 354 2390 594 2530
rect 974 2150 1005 2300
rect 1005 2150 1057 2300
rect 1057 2150 1201 2300
rect 1201 2150 1253 2300
rect 1253 2150 1374 2300
rect 984 1750 1005 1900
rect 1005 1750 1057 1900
rect 1057 1750 1201 1900
rect 1201 1750 1253 1900
rect 1253 1750 1384 1900
rect 354 1510 594 1650
rect 4660 1930 4740 2000
rect 2834 1653 3274 1670
rect 2834 1493 3047 1653
rect 3047 1493 3099 1653
rect 3099 1493 3274 1653
rect 2834 1490 3274 1493
rect 524 1078 844 1080
rect 524 918 533 1078
rect 533 918 677 1078
rect 677 918 729 1078
rect 729 918 844 1078
rect 524 910 844 918
rect 984 680 1023 830
rect 1023 680 1167 830
rect 1167 680 1219 830
rect 1219 680 1384 830
rect 2834 758 3274 770
rect 2834 598 2867 758
rect 2867 598 2919 758
rect 2919 598 3063 758
rect 3063 598 3115 758
rect 3115 598 3259 758
rect 3259 598 3274 758
rect 2834 590 3274 598
rect 984 310 1023 460
rect 1023 310 1167 460
rect 1167 310 1219 460
rect 1219 310 1384 460
rect 524 60 533 220
rect 533 60 677 220
rect 677 60 729 220
rect 729 60 844 220
rect 524 -366 844 60
rect 2834 -100 3274 -90
rect 2834 -260 2867 -100
rect 2867 -260 2919 -100
rect 2919 -260 3063 -100
rect 3063 -260 3115 -100
rect 3115 -260 3259 -100
rect 3259 -260 3274 -100
rect 2834 -270 3274 -260
rect 524 -526 533 -366
rect 533 -526 677 -366
rect 677 -526 729 -366
rect 729 -526 844 -366
rect 524 -530 844 -526
rect 984 -760 1023 -610
rect 1023 -760 1167 -610
rect 1167 -760 1219 -610
rect 1219 -760 1384 -610
rect 984 -984 1384 -980
rect 984 -1130 1023 -984
rect 1023 -1130 1167 -984
rect 1167 -1130 1219 -984
rect 1219 -1130 1384 -984
rect 524 -1224 844 -1220
rect 524 -1384 533 -1224
rect 533 -1384 677 -1224
rect 677 -1384 729 -1224
rect 729 -1384 844 -1224
rect 524 -1390 844 -1384
rect -146 -1786 174 -1770
rect -146 -1946 -97 -1786
rect -97 -1946 43 -1786
rect 43 -1946 95 -1786
rect 95 -1946 174 -1786
rect 3140 -1780 3320 -1660
rect -146 -1950 174 -1946
rect 524 -2186 575 -2030
rect 575 -2186 715 -2030
rect 715 -2186 767 -2030
rect 767 -2186 844 -2030
rect 524 -2404 844 -2186
rect 524 -2564 575 -2404
rect 575 -2564 715 -2404
rect 715 -2564 767 -2404
rect 767 -2564 844 -2404
rect 524 -2570 844 -2564
rect 1260 -2250 1344 -2150
rect 1344 -2250 1474 -2150
rect 1474 -2250 1530 -2150
rect 1260 -2420 1530 -2250
rect -146 -2804 -97 -2650
rect -97 -2804 43 -2650
rect 43 -2804 95 -2650
rect 95 -2804 174 -2650
rect -146 -3022 174 -2804
rect -146 -3182 -97 -3022
rect -97 -3182 43 -3022
rect 43 -3182 95 -3022
rect 95 -3182 174 -3022
rect -146 -3190 174 -3182
rect 524 -3262 844 -3260
rect 524 -3422 575 -3262
rect 575 -3422 715 -3262
rect 715 -3422 767 -3262
rect 767 -3422 844 -3262
rect 524 -3640 844 -3422
rect 524 -3800 575 -3640
rect 575 -3800 715 -3640
rect 715 -3800 767 -3640
rect 767 -3800 844 -3640
rect -146 -3880 174 -3870
rect -146 -4040 -97 -3880
rect -97 -4040 43 -3880
rect 43 -4040 95 -3880
rect 95 -4040 174 -3880
rect -146 -4050 174 -4040
rect 354 -4680 594 -4540
rect 974 -4920 1005 -4770
rect 1005 -4920 1057 -4770
rect 1057 -4920 1201 -4770
rect 1201 -4920 1253 -4770
rect 1253 -4920 1374 -4770
rect 984 -5320 1005 -5170
rect 1005 -5320 1057 -5170
rect 1057 -5320 1201 -5170
rect 1201 -5320 1253 -5170
rect 1253 -5320 1384 -5170
rect 354 -5560 594 -5420
rect 5080 -5200 5170 -5080
rect 2834 -5417 3274 -5400
rect 2834 -5577 3047 -5417
rect 3047 -5577 3099 -5417
rect 3099 -5577 3274 -5417
rect 2834 -5580 3274 -5577
rect 524 -5992 844 -5990
rect 524 -6152 533 -5992
rect 533 -6152 677 -5992
rect 677 -6152 729 -5992
rect 729 -6152 844 -5992
rect 524 -6160 844 -6152
rect 984 -6390 1023 -6240
rect 1023 -6390 1167 -6240
rect 1167 -6390 1219 -6240
rect 1219 -6390 1384 -6240
rect 2834 -6312 3274 -6300
rect 2834 -6472 2867 -6312
rect 2867 -6472 2919 -6312
rect 2919 -6472 3063 -6312
rect 3063 -6472 3115 -6312
rect 3115 -6472 3259 -6312
rect 3259 -6472 3274 -6312
rect 2834 -6480 3274 -6472
rect 984 -6760 1023 -6610
rect 1023 -6760 1167 -6610
rect 1167 -6760 1219 -6610
rect 1219 -6760 1384 -6610
rect 524 -7010 533 -6850
rect 533 -7010 677 -6850
rect 677 -7010 729 -6850
rect 729 -7010 844 -6850
rect 524 -7436 844 -7010
rect 2834 -7170 3274 -7160
rect 2834 -7330 2867 -7170
rect 2867 -7330 2919 -7170
rect 2919 -7330 3063 -7170
rect 3063 -7330 3115 -7170
rect 3115 -7330 3259 -7170
rect 3259 -7330 3274 -7170
rect 2834 -7340 3274 -7330
rect 524 -7596 533 -7436
rect 533 -7596 677 -7436
rect 677 -7596 729 -7436
rect 729 -7596 844 -7436
rect 524 -7600 844 -7596
rect 984 -7830 1023 -7680
rect 1023 -7830 1167 -7680
rect 1167 -7830 1219 -7680
rect 1219 -7830 1384 -7680
rect 984 -8054 1384 -8050
rect 984 -8200 1023 -8054
rect 1023 -8200 1167 -8054
rect 1167 -8200 1219 -8054
rect 1219 -8200 1384 -8054
rect 2850 -8140 3020 -7990
rect 4550 -8250 4557 -8090
rect 4557 -8250 4609 -8090
rect 4609 -8250 4620 -8090
rect 524 -8294 844 -8290
rect 524 -8454 533 -8294
rect 533 -8454 677 -8294
rect 677 -8454 729 -8294
rect 729 -8454 844 -8294
rect 524 -8460 844 -8454
rect -146 -8856 174 -8840
rect -146 -9016 -97 -8856
rect -97 -9016 43 -8856
rect 43 -9016 95 -8856
rect 95 -9016 174 -8856
rect -146 -9020 174 -9016
rect 524 -9256 575 -9100
rect 575 -9256 715 -9100
rect 715 -9256 767 -9100
rect 767 -9256 844 -9100
rect 524 -9474 844 -9256
rect 524 -9634 575 -9474
rect 575 -9634 715 -9474
rect 715 -9634 767 -9474
rect 767 -9634 844 -9474
rect 524 -9640 844 -9634
rect 1250 -9320 1344 -9210
rect 1344 -9320 1474 -9210
rect 1474 -9320 1480 -9210
rect 1250 -9650 1480 -9320
rect 6060 -9410 6130 -9300
rect -146 -9874 -97 -9720
rect -97 -9874 43 -9720
rect 43 -9874 95 -9720
rect 95 -9874 174 -9720
rect -146 -10092 174 -9874
rect 6390 -10070 6460 -9960
rect -146 -10252 -97 -10092
rect -97 -10252 43 -10092
rect 43 -10252 95 -10092
rect 95 -10252 174 -10092
rect -146 -10260 174 -10252
rect 524 -10332 844 -10330
rect 524 -10492 575 -10332
rect 575 -10492 715 -10332
rect 715 -10492 767 -10332
rect 767 -10492 844 -10332
rect 524 -10710 844 -10492
rect 524 -10870 575 -10710
rect 575 -10870 715 -10710
rect 715 -10870 767 -10710
rect 767 -10870 844 -10710
rect -146 -10950 174 -10940
rect -146 -11110 -97 -10950
rect -97 -11110 43 -10950
rect 43 -11110 95 -10950
rect 95 -11110 174 -10950
rect -146 -11120 174 -11110
<< metal3 >>
rect 354 2540 594 2550
rect 314 2200 324 2540
rect 644 2200 654 2540
rect 974 2305 1394 2310
rect 964 2300 1394 2305
rect 354 2030 594 2200
rect 964 2150 974 2300
rect 1374 2150 1394 2300
rect 964 2145 1394 2150
rect 344 1870 604 2030
rect 974 1900 1394 2145
rect 4630 1910 4640 2020
rect 4760 1910 4770 2020
rect 354 1655 594 1870
rect 974 1750 984 1900
rect 1384 1750 1394 1900
rect 344 1650 604 1655
rect 344 1510 354 1650
rect 594 1510 604 1650
rect 344 1505 604 1510
rect 514 1080 854 1085
rect 514 910 524 1080
rect 844 910 854 1080
rect 514 905 854 910
rect 524 225 844 905
rect 974 830 1394 1750
rect 2824 1670 3284 1675
rect 2824 1490 2834 1670
rect 3274 1490 3284 1670
rect 2824 1485 3284 1490
rect 974 680 984 830
rect 1384 680 1394 830
rect 2834 775 3274 1485
rect 974 460 1394 680
rect 2824 770 3284 775
rect 2824 590 2834 770
rect 3274 590 3284 770
rect 2824 585 3284 590
rect 974 310 984 460
rect 1384 310 1394 460
rect 974 305 1394 310
rect 514 220 854 225
rect 514 -530 524 220
rect 844 -530 854 220
rect 514 -535 854 -530
rect 974 120 1384 305
rect 524 -1215 844 -535
rect 974 -610 1394 120
rect 2834 -85 3274 585
rect 2824 -90 3284 -85
rect 2824 -270 2834 -90
rect 3274 -270 3284 -90
rect 2824 -275 3284 -270
rect 974 -760 984 -610
rect 1384 -760 1394 -610
rect 974 -980 1394 -760
rect 974 -1130 984 -980
rect 1384 -1130 1394 -980
rect 974 -1150 1394 -1130
rect 514 -1220 854 -1215
rect 514 -1390 524 -1220
rect 844 -1390 854 -1220
rect 514 -1395 854 -1390
rect -156 -1770 184 -1765
rect -156 -1950 -146 -1770
rect 174 -1950 184 -1770
rect -156 -1955 184 -1950
rect -146 -2110 174 -1955
rect 524 -2025 844 -1395
rect 3130 -1660 3330 -1650
rect 3130 -1780 3140 -1660
rect 3320 -1780 3330 -1660
rect 3130 -1990 3330 -1780
rect 1630 -2018 4929 -1990
rect 514 -2030 854 -2025
rect -156 -2260 184 -2110
rect 514 -2120 524 -2030
rect -156 -2570 -146 -2260
rect 174 -2570 184 -2260
rect 504 -2550 524 -2120
rect 514 -2570 524 -2550
rect 844 -2570 854 -2030
rect 1250 -2150 1540 -2145
rect 1250 -2420 1260 -2150
rect 1530 -2420 1540 -2150
rect 1250 -2425 1540 -2420
rect -146 -2645 174 -2570
rect 514 -2575 854 -2570
rect -156 -2650 184 -2645
rect -156 -3190 -146 -2650
rect 174 -3190 184 -2650
rect -156 -3195 184 -3190
rect -146 -3865 174 -3195
rect 524 -3255 844 -2575
rect 514 -3260 854 -3255
rect 514 -3800 524 -3260
rect 844 -3800 854 -3260
rect 514 -3805 854 -3800
rect -156 -3870 184 -3865
rect -156 -4050 -146 -3870
rect 174 -4050 184 -3870
rect -156 -4055 184 -4050
rect 354 -4530 594 -4520
rect 314 -4870 324 -4530
rect 644 -4870 654 -4530
rect 1630 -4562 4845 -2018
rect 4909 -4562 4929 -2018
rect 1630 -4590 4929 -4562
rect 974 -4765 1394 -4760
rect 964 -4770 1394 -4765
rect 354 -5040 594 -4870
rect 964 -4920 974 -4770
rect 1374 -4920 1394 -4770
rect 964 -4925 1394 -4920
rect 344 -5200 604 -5040
rect 974 -5170 1394 -4925
rect 354 -5415 594 -5200
rect 974 -5320 984 -5170
rect 1384 -5320 1394 -5170
rect 5070 -5080 5180 -5075
rect 5070 -5200 5080 -5080
rect 5170 -5200 5180 -5080
rect 5070 -5205 5180 -5200
rect 344 -5420 604 -5415
rect 344 -5560 354 -5420
rect 594 -5560 604 -5420
rect 344 -5565 604 -5560
rect 514 -5990 854 -5985
rect 514 -6160 524 -5990
rect 844 -6160 854 -5990
rect 514 -6165 854 -6160
rect 524 -6845 844 -6165
rect 974 -6240 1394 -5320
rect 2824 -5400 3284 -5395
rect 2824 -5580 2834 -5400
rect 3274 -5580 3284 -5400
rect 2824 -5585 3284 -5580
rect 974 -6390 984 -6240
rect 1384 -6390 1394 -6240
rect 2834 -6295 3274 -5585
rect 974 -6610 1394 -6390
rect 2824 -6300 3284 -6295
rect 2824 -6480 2834 -6300
rect 3274 -6480 3284 -6300
rect 2824 -6485 3284 -6480
rect 974 -6760 984 -6610
rect 1384 -6760 1394 -6610
rect 974 -6765 1394 -6760
rect 514 -6850 854 -6845
rect 514 -7600 524 -6850
rect 844 -7600 854 -6850
rect 514 -7605 854 -7600
rect 974 -6950 1384 -6765
rect 524 -8285 844 -7605
rect 974 -7680 1394 -6950
rect 2834 -7155 3274 -6485
rect 2824 -7160 3284 -7155
rect 2824 -7340 2834 -7160
rect 3274 -7340 3284 -7160
rect 2824 -7345 3284 -7340
rect 974 -7830 984 -7680
rect 1384 -7830 1394 -7680
rect 974 -8050 1394 -7830
rect 974 -8200 984 -8050
rect 1384 -8200 1394 -8050
rect 2840 -7990 3030 -7985
rect 2840 -8140 2850 -7990
rect 3020 -8140 3030 -7990
rect 2840 -8145 3030 -8140
rect 4540 -8090 4630 -8085
rect 974 -8220 1394 -8200
rect 514 -8290 854 -8285
rect 514 -8460 524 -8290
rect 844 -8460 854 -8290
rect 514 -8465 854 -8460
rect -156 -8840 184 -8835
rect -156 -9020 -146 -8840
rect 174 -9020 184 -8840
rect -156 -9025 184 -9020
rect -146 -9180 174 -9025
rect 524 -9095 844 -8465
rect 2850 -9080 3020 -8145
rect 4540 -8250 4550 -8090
rect 4620 -8250 5190 -8090
rect 4540 -8255 4630 -8250
rect 514 -9100 854 -9095
rect -156 -9330 184 -9180
rect 514 -9190 524 -9100
rect -156 -9640 -146 -9330
rect 174 -9640 184 -9330
rect 504 -9620 524 -9190
rect 514 -9640 524 -9620
rect 844 -9640 854 -9100
rect 1640 -9108 4939 -9080
rect -146 -9715 174 -9640
rect 514 -9645 854 -9640
rect 1240 -9210 1490 -9205
rect -156 -9720 184 -9715
rect -156 -10260 -146 -9720
rect 174 -10260 184 -9720
rect -156 -10265 184 -10260
rect -146 -10935 174 -10265
rect 524 -10325 844 -9645
rect 1240 -9650 1250 -9210
rect 1480 -9650 1490 -9210
rect 1240 -9655 1490 -9650
rect 514 -10330 854 -10325
rect 514 -10870 524 -10330
rect 844 -10870 854 -10330
rect 514 -10875 854 -10870
rect -156 -10940 184 -10935
rect -156 -11120 -146 -10940
rect 174 -11120 184 -10940
rect -156 -11125 184 -11120
rect 1640 -11652 4855 -9108
rect 4919 -11652 4939 -9108
rect 6050 -9300 6140 -9295
rect 6050 -9410 6060 -9300
rect 6130 -9410 6460 -9300
rect 6050 -9415 6140 -9410
rect 6390 -9955 6460 -9410
rect 6380 -9960 6470 -9955
rect 6380 -10070 6390 -9960
rect 6460 -10070 6470 -9960
rect 6380 -10075 6470 -10070
rect 1640 -11680 4939 -11652
<< via3 >>
rect 324 2530 644 2540
rect 324 2390 354 2530
rect 354 2390 594 2530
rect 594 2390 644 2530
rect 324 2200 644 2390
rect 4640 2000 4760 2020
rect 4640 1930 4660 2000
rect 4660 1930 4740 2000
rect 4740 1930 4760 2000
rect 4640 1910 4760 1930
rect -146 -2570 174 -2260
rect 1260 -2420 1530 -2150
rect 324 -4540 644 -4530
rect 324 -4680 354 -4540
rect 354 -4680 594 -4540
rect 594 -4680 644 -4540
rect 324 -4870 644 -4680
rect 4845 -4562 4909 -2018
rect 5080 -5200 5170 -5080
rect -146 -9640 174 -9330
rect 1250 -9650 1480 -9210
rect 4855 -11652 4919 -9108
<< mimcap >>
rect 1730 -2130 4730 -2090
rect 1730 -4450 1770 -2130
rect 4690 -4450 4730 -2130
rect 1730 -4490 4730 -4450
rect 1740 -9220 4740 -9180
rect 1740 -11540 1780 -9220
rect 4700 -11540 4740 -9220
rect 1740 -11580 4740 -11540
<< mimcapcontact >>
rect 1770 -4450 4690 -2130
rect 1780 -11540 4700 -9220
<< metal4 >>
rect 323 2540 645 2541
rect 323 2200 324 2540
rect 644 2200 645 2540
rect 323 2199 645 2200
rect 4639 2020 4761 2021
rect 4639 1910 4640 2020
rect 4760 1960 4761 2020
rect 5022 1960 11724 2001
rect 4760 1910 5042 1960
rect 4639 1909 5042 1910
rect 4640 1850 5042 1909
rect -1346 1729 4356 1770
rect -1346 -1989 4100 1729
rect 4336 -1989 4356 1729
rect -1346 -2030 4356 -1989
rect 4829 -2018 4925 -2002
rect 1769 -2130 4691 -2129
rect 1259 -2150 1531 -2149
rect -147 -2260 175 -2259
rect 1259 -2260 1260 -2150
rect 1530 -2260 1531 -2150
rect 1769 -2260 1770 -2130
rect -147 -2570 -146 -2260
rect 174 -2570 175 -2260
rect 1530 -2420 1770 -2260
rect 1370 -2560 1770 -2420
rect -147 -2571 175 -2570
rect 1769 -4450 1770 -2560
rect 4690 -4450 4691 -2130
rect 1769 -4451 4691 -4450
rect 323 -4530 645 -4529
rect 323 -4870 324 -4530
rect 644 -4870 645 -4530
rect 4829 -4562 4845 -2018
rect 4909 -4562 4925 -2018
rect 5022 -4158 5042 1850
rect 5278 -4158 11724 1960
rect 5022 -4190 11724 -4158
rect 5022 -4199 11730 -4190
rect 4829 -4578 4925 -4562
rect 323 -4871 645 -4870
rect 5060 -5080 5760 -4199
rect 5060 -5200 5080 -5080
rect 5170 -5200 5760 -5080
rect -1346 -5341 4356 -5300
rect 5060 -5309 5760 -5200
rect 11390 -5309 11730 -4199
rect -1346 -9059 4100 -5341
rect 4336 -9059 4356 -5341
rect -1346 -9100 4356 -9059
rect 5022 -5310 11730 -5309
rect 5022 -5350 11724 -5310
rect 4839 -9108 4935 -9092
rect 1249 -9210 1481 -9209
rect -147 -9330 175 -9329
rect -147 -9640 -146 -9330
rect 174 -9640 175 -9330
rect 1249 -9380 1250 -9210
rect 1480 -9380 1481 -9210
rect 1779 -9220 4701 -9219
rect 1779 -9380 1780 -9220
rect -147 -9641 175 -9640
rect 1480 -9650 1780 -9380
rect 1360 -9800 1780 -9650
rect 1779 -11540 1780 -9800
rect 4700 -11540 4701 -9220
rect 1779 -11541 4701 -11540
rect 4839 -11652 4855 -9108
rect 4919 -11652 4935 -9108
rect 5022 -11468 5042 -5350
rect 5278 -11468 11724 -5350
rect 5022 -11509 11724 -11468
rect 4839 -11668 4935 -11652
<< via4 >>
rect 324 2200 644 2540
rect 4100 -1989 4336 1729
rect -146 -2570 174 -2260
rect 1090 -2420 1260 -2260
rect 1260 -2420 1370 -2260
rect 1090 -2560 1370 -2420
rect 324 -4870 644 -4530
rect 5042 -4158 5278 1960
rect 4100 -9059 4336 -5341
rect -146 -9640 174 -9330
rect 1060 -9650 1250 -9380
rect 1250 -9650 1360 -9380
rect 1060 -9800 1360 -9650
rect 5042 -11468 5278 -5350
<< mimcap2 >>
rect 5624 1861 11624 1901
rect -1246 1630 3754 1670
rect -1246 -1890 -1206 1630
rect 3714 -1890 3754 1630
rect -1246 -1930 3754 -1890
rect 5624 -4059 5664 1861
rect 11584 -4059 11624 1861
rect 5624 -4099 11624 -4059
rect -1246 -5440 3754 -5400
rect -1246 -8960 -1206 -5440
rect 3714 -8960 3754 -5440
rect -1246 -9000 3754 -8960
rect 5624 -5449 11624 -5409
rect 5624 -11369 5664 -5449
rect 11584 -11369 11624 -5449
rect 5624 -11409 11624 -11369
<< mimcap2contact >>
rect -1206 -1890 3714 1630
rect 5664 -4059 11584 1861
rect -1206 -8960 3714 -5440
rect 5664 -11369 11584 -5449
<< metal5 >>
rect 294 2540 674 2570
rect 294 2200 324 2540
rect 644 2200 674 2540
rect 294 1654 674 2200
rect 3230 2360 5960 2680
rect 3230 1654 3590 2360
rect 5000 1960 5320 2002
rect 4058 1729 4378 1771
rect -1230 1630 3738 1654
rect -1230 -1890 -1206 1630
rect 3714 -1890 3738 1630
rect -1230 -1914 3738 -1890
rect 4058 -1989 4100 1729
rect 4336 -1989 4378 1729
rect 4058 -2031 4378 -1989
rect -170 -2240 198 -2236
rect 1066 -2240 1394 -2236
rect -170 -2260 3564 -2240
rect -170 -2570 -146 -2260
rect 174 -2560 1090 -2260
rect 1370 -2360 3564 -2260
rect 5000 -2360 5042 1960
rect 1370 -2560 5042 -2360
rect 174 -2570 198 -2560
rect -170 -2594 198 -2570
rect 1066 -2584 1394 -2560
rect 3224 -2680 5042 -2560
rect 5000 -4158 5042 -2680
rect 5278 -4158 5320 1960
rect 5640 1885 5960 2360
rect 5640 1861 11608 1885
rect 5640 -4059 5664 1861
rect 11584 -4059 11608 1861
rect 5640 -4083 11608 -4059
rect 5000 -4200 5320 -4158
rect 294 -4530 674 -4500
rect 294 -4870 324 -4530
rect 644 -4870 674 -4530
rect 5750 -4590 6070 -4083
rect 294 -5416 674 -4870
rect 3300 -4970 6070 -4590
rect 3300 -5416 3680 -4970
rect 4680 -4980 6070 -4970
rect 4058 -5341 4378 -5299
rect -1230 -5440 3738 -5416
rect -1230 -8960 -1206 -5440
rect 3714 -8960 3738 -5440
rect -1230 -8984 3738 -8960
rect 4058 -9059 4100 -5341
rect 4336 -9059 4378 -5341
rect 4058 -9101 4378 -9059
rect 5000 -5350 5320 -5308
rect -170 -9310 198 -9306
rect -170 -9330 3564 -9310
rect -170 -9640 -146 -9330
rect 174 -9380 3564 -9330
rect 174 -9630 1060 -9380
rect 174 -9640 198 -9630
rect -170 -9664 198 -9640
rect 1036 -9800 1060 -9630
rect 1360 -9430 3564 -9380
rect 5000 -9430 5042 -5350
rect 1360 -9630 5042 -9430
rect 1360 -9800 1384 -9630
rect 3224 -9750 5042 -9630
rect 1036 -9824 1384 -9800
rect 5000 -11468 5042 -9750
rect 5278 -11468 5320 -5350
rect 5750 -5425 6070 -4980
rect 11110 -5425 11470 -4083
rect 5640 -5449 11608 -5425
rect 5640 -11369 5664 -5449
rect 11584 -11369 11608 -5449
rect 5640 -11393 11608 -11369
rect 5000 -11510 5320 -11468
<< labels >>
rlabel metal1 -1840 -1240 -1560 -1040 1 Input
port 6 n
rlabel metal4 11480 -4560 11690 -4360 1 VN
port 8 n
rlabel metal2 2720 -1460 2890 -1320 3 VM5D
rlabel metal3 1040 1990 1140 2120 1 Out_1
port 4 n
rlabel metal2 4600 -8760 4720 -8660 1 VM6D
rlabel metal3 6390 -9510 6450 -9410 1 Disable_TIA
port 5 n
rlabel metal1 6090 -9890 6150 -9850 1 Disable_TIA_B
rlabel metal3 630 -10020 700 -9920 1 VM40D
rlabel metal3 630 -2970 700 -2870 1 VM28D
rlabel metal3 5080 -8250 5190 -8090 1 I_Bias1
port 7 n
rlabel metal2 1800 670 1910 840 1 Out_1
rlabel metal3 2900 1040 3170 1170 1 Out_2
port 2 n
rlabel metal5 11130 -5060 11230 -4890 1 VPP
port 1 n
<< end >>
