** sch_path: /home/simon/code/caravel_tia/xschem/test.sch
**.subckt test
x1 __UNCONNECTED_PIN__0 __UNCONNECTED_PIN__1 __UNCONNECTED_PIN__2 __UNCONNECTED_PIN__3
+ __UNCONNECTED_PIN__4 __UNCONNECTED_PIN__5 __UNCONNECTED_PIN__6 __UNCONNECTED_PIN__7 __UNCONNECTED_PIN__8
+ __UNCONNECTED_PIN__9 __UNCONNECTED_PIN__10 __UNCONNECTED_PIN__11 __UNCONNECTED_PIN__12 __UNCONNECTED_PIN__13[3]
+ __UNCONNECTED_PIN__13[2] __UNCONNECTED_PIN__13[1] __UNCONNECTED_PIN__13[0] __UNCONNECTED_PIN__14[31]
+ __UNCONNECTED_PIN__14[30] __UNCONNECTED_PIN__14[29] __UNCONNECTED_PIN__14[28] __UNCONNECTED_PIN__14[27]
+ __UNCONNECTED_PIN__14[26] __UNCONNECTED_PIN__14[25] __UNCONNECTED_PIN__14[24] __UNCONNECTED_PIN__14[23]
+ __UNCONNECTED_PIN__14[22] __UNCONNECTED_PIN__14[21] __UNCONNECTED_PIN__14[20] __UNCONNECTED_PIN__14[19]
+ __UNCONNECTED_PIN__14[18] __UNCONNECTED_PIN__14[17] __UNCONNECTED_PIN__14[16] __UNCONNECTED_PIN__14[15]
+ __UNCONNECTED_PIN__14[14] __UNCONNECTED_PIN__14[13] __UNCONNECTED_PIN__14[12] __UNCONNECTED_PIN__14[11]
+ __UNCONNECTED_PIN__14[10] __UNCONNECTED_PIN__14[9] __UNCONNECTED_PIN__14[8] __UNCONNECTED_PIN__14[7] __UNCONNECTED_PIN__14[6]
+ __UNCONNECTED_PIN__14[5] __UNCONNECTED_PIN__14[4] __UNCONNECTED_PIN__14[3] __UNCONNECTED_PIN__14[2] __UNCONNECTED_PIN__14[1]
+ __UNCONNECTED_PIN__14[0] __UNCONNECTED_PIN__15[31] __UNCONNECTED_PIN__15[30] __UNCONNECTED_PIN__15[29]
+ __UNCONNECTED_PIN__15[28] __UNCONNECTED_PIN__15[27] __UNCONNECTED_PIN__15[26] __UNCONNECTED_PIN__15[25]
+ __UNCONNECTED_PIN__15[24] __UNCONNECTED_PIN__15[23] __UNCONNECTED_PIN__15[22] __UNCONNECTED_PIN__15[21]
+ __UNCONNECTED_PIN__15[20] __UNCONNECTED_PIN__15[19] __UNCONNECTED_PIN__15[18] __UNCONNECTED_PIN__15[17]
+ __UNCONNECTED_PIN__15[16] __UNCONNECTED_PIN__15[15] __UNCONNECTED_PIN__15[14] __UNCONNECTED_PIN__15[13]
+ __UNCONNECTED_PIN__15[12] __UNCONNECTED_PIN__15[11] __UNCONNECTED_PIN__15[10] __UNCONNECTED_PIN__15[9]
+ __UNCONNECTED_PIN__15[8] __UNCONNECTED_PIN__15[7] __UNCONNECTED_PIN__15[6] __UNCONNECTED_PIN__15[5] __UNCONNECTED_PIN__15[4]
+ __UNCONNECTED_PIN__15[3] __UNCONNECTED_PIN__15[2] __UNCONNECTED_PIN__15[1] __UNCONNECTED_PIN__15[0] __UNCONNECTED_PIN__16
+ __UNCONNECTED_PIN__17[31] __UNCONNECTED_PIN__17[30] __UNCONNECTED_PIN__17[29] __UNCONNECTED_PIN__17[28]
+ __UNCONNECTED_PIN__17[27] __UNCONNECTED_PIN__17[26] __UNCONNECTED_PIN__17[25] __UNCONNECTED_PIN__17[24]
+ __UNCONNECTED_PIN__17[23] __UNCONNECTED_PIN__17[22] __UNCONNECTED_PIN__17[21] __UNCONNECTED_PIN__17[20]
+ __UNCONNECTED_PIN__17[19] __UNCONNECTED_PIN__17[18] __UNCONNECTED_PIN__17[17] __UNCONNECTED_PIN__17[16]
+ __UNCONNECTED_PIN__17[15] __UNCONNECTED_PIN__17[14] __UNCONNECTED_PIN__17[13] __UNCONNECTED_PIN__17[12]
+ __UNCONNECTED_PIN__17[11] __UNCONNECTED_PIN__17[10] __UNCONNECTED_PIN__17[9] __UNCONNECTED_PIN__17[8]
+ __UNCONNECTED_PIN__17[7] __UNCONNECTED_PIN__17[6] __UNCONNECTED_PIN__17[5] __UNCONNECTED_PIN__17[4] __UNCONNECTED_PIN__17[3]
+ __UNCONNECTED_PIN__17[2] __UNCONNECTED_PIN__17[1] __UNCONNECTED_PIN__17[0] __UNCONNECTED_PIN__18[127]
+ __UNCONNECTED_PIN__18[126] __UNCONNECTED_PIN__18[125] __UNCONNECTED_PIN__18[124] __UNCONNECTED_PIN__18[123]
+ __UNCONNECTED_PIN__18[122] __UNCONNECTED_PIN__18[121] __UNCONNECTED_PIN__18[120] __UNCONNECTED_PIN__18[119]
+ __UNCONNECTED_PIN__18[118] __UNCONNECTED_PIN__18[117] __UNCONNECTED_PIN__18[116] __UNCONNECTED_PIN__18[115]
+ __UNCONNECTED_PIN__18[114] __UNCONNECTED_PIN__18[113] __UNCONNECTED_PIN__18[112] __UNCONNECTED_PIN__18[111]
+ __UNCONNECTED_PIN__18[110] __UNCONNECTED_PIN__18[109] __UNCONNECTED_PIN__18[108] __UNCONNECTED_PIN__18[107]
+ __UNCONNECTED_PIN__18[106] __UNCONNECTED_PIN__18[105] __UNCONNECTED_PIN__18[104] __UNCONNECTED_PIN__18[103]
+ __UNCONNECTED_PIN__18[102] __UNCONNECTED_PIN__18[101] __UNCONNECTED_PIN__18[100] __UNCONNECTED_PIN__18[99]
+ __UNCONNECTED_PIN__18[98] __UNCONNECTED_PIN__18[97] __UNCONNECTED_PIN__18[96] __UNCONNECTED_PIN__18[95]
+ __UNCONNECTED_PIN__18[94] __UNCONNECTED_PIN__18[93] __UNCONNECTED_PIN__18[92] __UNCONNECTED_PIN__18[91]
+ __UNCONNECTED_PIN__18[90] __UNCONNECTED_PIN__18[89] __UNCONNECTED_PIN__18[88] __UNCONNECTED_PIN__18[87]
+ __UNCONNECTED_PIN__18[86] __UNCONNECTED_PIN__18[85] __UNCONNECTED_PIN__18[84] __UNCONNECTED_PIN__18[83]
+ __UNCONNECTED_PIN__18[82] __UNCONNECTED_PIN__18[81] __UNCONNECTED_PIN__18[80] __UNCONNECTED_PIN__18[79]
+ __UNCONNECTED_PIN__18[78] __UNCONNECTED_PIN__18[77] __UNCONNECTED_PIN__18[76] __UNCONNECTED_PIN__18[75]
+ __UNCONNECTED_PIN__18[74] __UNCONNECTED_PIN__18[73] __UNCONNECTED_PIN__18[72] __UNCONNECTED_PIN__18[71]
+ __UNCONNECTED_PIN__18[70] __UNCONNECTED_PIN__18[69] __UNCONNECTED_PIN__18[68] __UNCONNECTED_PIN__18[67]
+ __UNCONNECTED_PIN__18[66] __UNCONNECTED_PIN__18[65] __UNCONNECTED_PIN__18[64] __UNCONNECTED_PIN__18[63]
+ __UNCONNECTED_PIN__18[62] __UNCONNECTED_PIN__18[61] __UNCONNECTED_PIN__18[60] __UNCONNECTED_PIN__18[59]
+ __UNCONNECTED_PIN__18[58] __UNCONNECTED_PIN__18[57] __UNCONNECTED_PIN__18[56] __UNCONNECTED_PIN__18[55]
+ __UNCONNECTED_PIN__18[54] __UNCONNECTED_PIN__18[53] __UNCONNECTED_PIN__18[52] __UNCONNECTED_PIN__18[51]
+ __UNCONNECTED_PIN__18[50] __UNCONNECTED_PIN__18[49] __UNCONNECTED_PIN__18[48] __UNCONNECTED_PIN__18[47]
+ __UNCONNECTED_PIN__18[46] __UNCONNECTED_PIN__18[45] __UNCONNECTED_PIN__18[44] __UNCONNECTED_PIN__18[43]
+ __UNCONNECTED_PIN__18[42] __UNCONNECTED_PIN__18[41] __UNCONNECTED_PIN__18[40] __UNCONNECTED_PIN__18[39]
+ __UNCONNECTED_PIN__18[38] __UNCONNECTED_PIN__18[37] __UNCONNECTED_PIN__18[36] __UNCONNECTED_PIN__18[35]
+ __UNCONNECTED_PIN__18[34] __UNCONNECTED_PIN__18[33] __UNCONNECTED_PIN__18[32] __UNCONNECTED_PIN__18[31]
+ __UNCONNECTED_PIN__18[30] __UNCONNECTED_PIN__18[29] __UNCONNECTED_PIN__18[28] __UNCONNECTED_PIN__18[27]
+ __UNCONNECTED_PIN__18[26] __UNCONNECTED_PIN__18[25] __UNCONNECTED_PIN__18[24] __UNCONNECTED_PIN__18[23]
+ __UNCONNECTED_PIN__18[22] __UNCONNECTED_PIN__18[21] __UNCONNECTED_PIN__18[20] __UNCONNECTED_PIN__18[19]
+ __UNCONNECTED_PIN__18[18] __UNCONNECTED_PIN__18[17] __UNCONNECTED_PIN__18[16] __UNCONNECTED_PIN__18[15]
+ __UNCONNECTED_PIN__18[14] __UNCONNECTED_PIN__18[13] __UNCONNECTED_PIN__18[12] __UNCONNECTED_PIN__18[11]
+ __UNCONNECTED_PIN__18[10] __UNCONNECTED_PIN__18[9] __UNCONNECTED_PIN__18[8] __UNCONNECTED_PIN__18[7] __UNCONNECTED_PIN__18[6]
+ __UNCONNECTED_PIN__18[5] __UNCONNECTED_PIN__18[4] __UNCONNECTED_PIN__18[3] __UNCONNECTED_PIN__18[2] __UNCONNECTED_PIN__18[1]
+ __UNCONNECTED_PIN__18[0] __UNCONNECTED_PIN__19[127] __UNCONNECTED_PIN__19[126] __UNCONNECTED_PIN__19[125]
+ __UNCONNECTED_PIN__19[124] __UNCONNECTED_PIN__19[123] __UNCONNECTED_PIN__19[122] __UNCONNECTED_PIN__19[121]
+ __UNCONNECTED_PIN__19[120] __UNCONNECTED_PIN__19[119] __UNCONNECTED_PIN__19[118] __UNCONNECTED_PIN__19[117]
+ __UNCONNECTED_PIN__19[116] __UNCONNECTED_PIN__19[115] __UNCONNECTED_PIN__19[114] __UNCONNECTED_PIN__19[113]
+ __UNCONNECTED_PIN__19[112] __UNCONNECTED_PIN__19[111] __UNCONNECTED_PIN__19[110] __UNCONNECTED_PIN__19[109]
+ __UNCONNECTED_PIN__19[108] __UNCONNECTED_PIN__19[107] __UNCONNECTED_PIN__19[106] __UNCONNECTED_PIN__19[105]
+ __UNCONNECTED_PIN__19[104] __UNCONNECTED_PIN__19[103] __UNCONNECTED_PIN__19[102] __UNCONNECTED_PIN__19[101]
+ __UNCONNECTED_PIN__19[100] __UNCONNECTED_PIN__19[99] __UNCONNECTED_PIN__19[98] __UNCONNECTED_PIN__19[97]
+ __UNCONNECTED_PIN__19[96] __UNCONNECTED_PIN__19[95] __UNCONNECTED_PIN__19[94] __UNCONNECTED_PIN__19[93]
+ __UNCONNECTED_PIN__19[92] __UNCONNECTED_PIN__19[91] __UNCONNECTED_PIN__19[90] __UNCONNECTED_PIN__19[89]
+ __UNCONNECTED_PIN__19[88] __UNCONNECTED_PIN__19[87] __UNCONNECTED_PIN__19[86] __UNCONNECTED_PIN__19[85]
+ __UNCONNECTED_PIN__19[84] __UNCONNECTED_PIN__19[83] __UNCONNECTED_PIN__19[82] __UNCONNECTED_PIN__19[81]
+ __UNCONNECTED_PIN__19[80] __UNCONNECTED_PIN__19[79] __UNCONNECTED_PIN__19[78] __UNCONNECTED_PIN__19[77]
+ __UNCONNECTED_PIN__19[76] __UNCONNECTED_PIN__19[75] __UNCONNECTED_PIN__19[74] __UNCONNECTED_PIN__19[73]
+ __UNCONNECTED_PIN__19[72] __UNCONNECTED_PIN__19[71] __UNCONNECTED_PIN__19[70] __UNCONNECTED_PIN__19[69]
+ __UNCONNECTED_PIN__19[68] __UNCONNECTED_PIN__19[67] __UNCONNECTED_PIN__19[66] __UNCONNECTED_PIN__19[65]
+ __UNCONNECTED_PIN__19[64] __UNCONNECTED_PIN__19[63] __UNCONNECTED_PIN__19[62] __UNCONNECTED_PIN__19[61]
+ __UNCONNECTED_PIN__19[60] __UNCONNECTED_PIN__19[59] __UNCONNECTED_PIN__19[58] __UNCONNECTED_PIN__19[57]
+ __UNCONNECTED_PIN__19[56] __UNCONNECTED_PIN__19[55] __UNCONNECTED_PIN__19[54] __UNCONNECTED_PIN__19[53]
+ __UNCONNECTED_PIN__19[52] __UNCONNECTED_PIN__19[51] __UNCONNECTED_PIN__19[50] __UNCONNECTED_PIN__19[49]
+ __UNCONNECTED_PIN__19[48] __UNCONNECTED_PIN__19[47] __UNCONNECTED_PIN__19[46] __UNCONNECTED_PIN__19[45]
+ __UNCONNECTED_PIN__19[44] __UNCONNECTED_PIN__19[43] __UNCONNECTED_PIN__19[42] __UNCONNECTED_PIN__19[41]
+ __UNCONNECTED_PIN__19[40] __UNCONNECTED_PIN__19[39] __UNCONNECTED_PIN__19[38] __UNCONNECTED_PIN__19[37]
+ __UNCONNECTED_PIN__19[36] __UNCONNECTED_PIN__19[35] __UNCONNECTED_PIN__19[34] __UNCONNECTED_PIN__19[33]
+ __UNCONNECTED_PIN__19[32] __UNCONNECTED_PIN__19[31] __UNCONNECTED_PIN__19[30] __UNCONNECTED_PIN__19[29]
+ __UNCONNECTED_PIN__19[28] __UNCONNECTED_PIN__19[27] __UNCONNECTED_PIN__19[26] __UNCONNECTED_PIN__19[25]
+ __UNCONNECTED_PIN__19[24] __UNCONNECTED_PIN__19[23] __UNCONNECTED_PIN__19[22] __UNCONNECTED_PIN__19[21]
+ __UNCONNECTED_PIN__19[20] __UNCONNECTED_PIN__19[19] __UNCONNECTED_PIN__19[18] __UNCONNECTED_PIN__19[17]
+ __UNCONNECTED_PIN__19[16] __UNCONNECTED_PIN__19[15] __UNCONNECTED_PIN__19[14] __UNCONNECTED_PIN__19[13]
+ __UNCONNECTED_PIN__19[12] __UNCONNECTED_PIN__19[11] __UNCONNECTED_PIN__19[10] __UNCONNECTED_PIN__19[9]
+ __UNCONNECTED_PIN__19[8] __UNCONNECTED_PIN__19[7] __UNCONNECTED_PIN__19[6] __UNCONNECTED_PIN__19[5] __UNCONNECTED_PIN__19[4]
+ __UNCONNECTED_PIN__19[3] __UNCONNECTED_PIN__19[2] __UNCONNECTED_PIN__19[1] __UNCONNECTED_PIN__19[0]
+ __UNCONNECTED_PIN__20[127] __UNCONNECTED_PIN__20[126] __UNCONNECTED_PIN__20[125] __UNCONNECTED_PIN__20[124]
+ __UNCONNECTED_PIN__20[123] __UNCONNECTED_PIN__20[122] __UNCONNECTED_PIN__20[121] __UNCONNECTED_PIN__20[120]
+ __UNCONNECTED_PIN__20[119] __UNCONNECTED_PIN__20[118] __UNCONNECTED_PIN__20[117] __UNCONNECTED_PIN__20[116]
+ __UNCONNECTED_PIN__20[115] __UNCONNECTED_PIN__20[114] __UNCONNECTED_PIN__20[113] __UNCONNECTED_PIN__20[112]
+ __UNCONNECTED_PIN__20[111] __UNCONNECTED_PIN__20[110] __UNCONNECTED_PIN__20[109] __UNCONNECTED_PIN__20[108]
+ __UNCONNECTED_PIN__20[107] __UNCONNECTED_PIN__20[106] __UNCONNECTED_PIN__20[105] __UNCONNECTED_PIN__20[104]
+ __UNCONNECTED_PIN__20[103] __UNCONNECTED_PIN__20[102] __UNCONNECTED_PIN__20[101] __UNCONNECTED_PIN__20[100]
+ __UNCONNECTED_PIN__20[99] __UNCONNECTED_PIN__20[98] __UNCONNECTED_PIN__20[97] __UNCONNECTED_PIN__20[96]
+ __UNCONNECTED_PIN__20[95] __UNCONNECTED_PIN__20[94] __UNCONNECTED_PIN__20[93] __UNCONNECTED_PIN__20[92]
+ __UNCONNECTED_PIN__20[91] __UNCONNECTED_PIN__20[90] __UNCONNECTED_PIN__20[89] __UNCONNECTED_PIN__20[88]
+ __UNCONNECTED_PIN__20[87] __UNCONNECTED_PIN__20[86] __UNCONNECTED_PIN__20[85] __UNCONNECTED_PIN__20[84]
+ __UNCONNECTED_PIN__20[83] __UNCONNECTED_PIN__20[82] __UNCONNECTED_PIN__20[81] __UNCONNECTED_PIN__20[80]
+ __UNCONNECTED_PIN__20[79] __UNCONNECTED_PIN__20[78] __UNCONNECTED_PIN__20[77] __UNCONNECTED_PIN__20[76]
+ __UNCONNECTED_PIN__20[75] __UNCONNECTED_PIN__20[74] __UNCONNECTED_PIN__20[73] __UNCONNECTED_PIN__20[72]
+ __UNCONNECTED_PIN__20[71] __UNCONNECTED_PIN__20[70] __UNCONNECTED_PIN__20[69] __UNCONNECTED_PIN__20[68]
+ __UNCONNECTED_PIN__20[67] __UNCONNECTED_PIN__20[66] __UNCONNECTED_PIN__20[65] __UNCONNECTED_PIN__20[64]
+ __UNCONNECTED_PIN__20[63] __UNCONNECTED_PIN__20[62] __UNCONNECTED_PIN__20[61] __UNCONNECTED_PIN__20[60]
+ __UNCONNECTED_PIN__20[59] __UNCONNECTED_PIN__20[58] __UNCONNECTED_PIN__20[57] __UNCONNECTED_PIN__20[56]
+ __UNCONNECTED_PIN__20[55] __UNCONNECTED_PIN__20[54] __UNCONNECTED_PIN__20[53] __UNCONNECTED_PIN__20[52]
+ __UNCONNECTED_PIN__20[51] __UNCONNECTED_PIN__20[50] __UNCONNECTED_PIN__20[49] __UNCONNECTED_PIN__20[48]
+ __UNCONNECTED_PIN__20[47] __UNCONNECTED_PIN__20[46] __UNCONNECTED_PIN__20[45] __UNCONNECTED_PIN__20[44]
+ __UNCONNECTED_PIN__20[43] __UNCONNECTED_PIN__20[42] __UNCONNECTED_PIN__20[41] __UNCONNECTED_PIN__20[40]
+ __UNCONNECTED_PIN__20[39] __UNCONNECTED_PIN__20[38] __UNCONNECTED_PIN__20[37] __UNCONNECTED_PIN__20[36]
+ __UNCONNECTED_PIN__20[35] __UNCONNECTED_PIN__20[34] __UNCONNECTED_PIN__20[33] __UNCONNECTED_PIN__20[32]
+ __UNCONNECTED_PIN__20[31] __UNCONNECTED_PIN__20[30] __UNCONNECTED_PIN__20[29] __UNCONNECTED_PIN__20[28]
+ __UNCONNECTED_PIN__20[27] __UNCONNECTED_PIN__20[26] __UNCONNECTED_PIN__20[25] __UNCONNECTED_PIN__20[24]
+ __UNCONNECTED_PIN__20[23] __UNCONNECTED_PIN__20[22] __UNCONNECTED_PIN__20[21] __UNCONNECTED_PIN__20[20]
+ __UNCONNECTED_PIN__20[19] __UNCONNECTED_PIN__20[18] __UNCONNECTED_PIN__20[17] __UNCONNECTED_PIN__20[16]
+ __UNCONNECTED_PIN__20[15] __UNCONNECTED_PIN__20[14] __UNCONNECTED_PIN__20[13] __UNCONNECTED_PIN__20[12]
+ __UNCONNECTED_PIN__20[11] __UNCONNECTED_PIN__20[10] __UNCONNECTED_PIN__20[9] __UNCONNECTED_PIN__20[8]
+ __UNCONNECTED_PIN__20[7] __UNCONNECTED_PIN__20[6] __UNCONNECTED_PIN__20[5] __UNCONNECTED_PIN__20[4] __UNCONNECTED_PIN__20[3]
+ __UNCONNECTED_PIN__20[2] __UNCONNECTED_PIN__20[1] __UNCONNECTED_PIN__20[0] __UNCONNECTED_PIN__21[26]
+ __UNCONNECTED_PIN__21[25] __UNCONNECTED_PIN__21[24] __UNCONNECTED_PIN__21[23] __UNCONNECTED_PIN__21[22]
+ __UNCONNECTED_PIN__21[21] __UNCONNECTED_PIN__21[20] __UNCONNECTED_PIN__21[19] __UNCONNECTED_PIN__21[18]
+ __UNCONNECTED_PIN__21[17] __UNCONNECTED_PIN__21[16] __UNCONNECTED_PIN__21[15] __UNCONNECTED_PIN__21[14]
+ __UNCONNECTED_PIN__21[13] __UNCONNECTED_PIN__21[12] __UNCONNECTED_PIN__21[11] __UNCONNECTED_PIN__21[10]
+ __UNCONNECTED_PIN__21[9] __UNCONNECTED_PIN__21[8] __UNCONNECTED_PIN__21[7] __UNCONNECTED_PIN__21[6] __UNCONNECTED_PIN__21[5]
+ __UNCONNECTED_PIN__21[4] __UNCONNECTED_PIN__21[3] __UNCONNECTED_PIN__21[2] __UNCONNECTED_PIN__21[1] __UNCONNECTED_PIN__21[0]
+ __UNCONNECTED_PIN__22[26] __UNCONNECTED_PIN__22[25] __UNCONNECTED_PIN__22[24] __UNCONNECTED_PIN__22[23]
+ __UNCONNECTED_PIN__22[22] __UNCONNECTED_PIN__22[21] __UNCONNECTED_PIN__22[20] __UNCONNECTED_PIN__22[19]
+ __UNCONNECTED_PIN__22[18] __UNCONNECTED_PIN__22[17] __UNCONNECTED_PIN__22[16] __UNCONNECTED_PIN__22[15]
+ __UNCONNECTED_PIN__22[14] __UNCONNECTED_PIN__22[13] __UNCONNECTED_PIN__22[12] __UNCONNECTED_PIN__22[11]
+ __UNCONNECTED_PIN__22[10] __UNCONNECTED_PIN__22[9] __UNCONNECTED_PIN__22[8] __UNCONNECTED_PIN__22[7] __UNCONNECTED_PIN__22[6]
+ __UNCONNECTED_PIN__22[5] __UNCONNECTED_PIN__22[4] __UNCONNECTED_PIN__22[3] __UNCONNECTED_PIN__22[2] __UNCONNECTED_PIN__22[1]
+ __UNCONNECTED_PIN__22[0] __UNCONNECTED_PIN__23[26] __UNCONNECTED_PIN__23[25] __UNCONNECTED_PIN__23[24]
+ __UNCONNECTED_PIN__23[23] __UNCONNECTED_PIN__23[22] __UNCONNECTED_PIN__23[21] __UNCONNECTED_PIN__23[20]
+ __UNCONNECTED_PIN__23[19] __UNCONNECTED_PIN__23[18] __UNCONNECTED_PIN__23[17] __UNCONNECTED_PIN__23[16]
+ __UNCONNECTED_PIN__23[15] __UNCONNECTED_PIN__23[14] __UNCONNECTED_PIN__23[13] __UNCONNECTED_PIN__23[12]
+ __UNCONNECTED_PIN__23[11] __UNCONNECTED_PIN__23[10] __UNCONNECTED_PIN__23[9] __UNCONNECTED_PIN__23[8]
+ __UNCONNECTED_PIN__23[7] __UNCONNECTED_PIN__23[6] __UNCONNECTED_PIN__23[5] __UNCONNECTED_PIN__23[4] __UNCONNECTED_PIN__23[3]
+ __UNCONNECTED_PIN__23[2] __UNCONNECTED_PIN__23[1] __UNCONNECTED_PIN__23[0] __UNCONNECTED_PIN__24[26]
+ __UNCONNECTED_PIN__24[25] __UNCONNECTED_PIN__24[24] __UNCONNECTED_PIN__24[23] __UNCONNECTED_PIN__24[22]
+ __UNCONNECTED_PIN__24[21] __UNCONNECTED_PIN__24[20] __UNCONNECTED_PIN__24[19] __UNCONNECTED_PIN__24[18]
+ __UNCONNECTED_PIN__24[17] __UNCONNECTED_PIN__24[16] __UNCONNECTED_PIN__24[15] __UNCONNECTED_PIN__24[14]
+ __UNCONNECTED_PIN__24[13] __UNCONNECTED_PIN__24[12] __UNCONNECTED_PIN__24[11] __UNCONNECTED_PIN__24[10]
+ __UNCONNECTED_PIN__24[9] __UNCONNECTED_PIN__24[8] __UNCONNECTED_PIN__24[7] __UNCONNECTED_PIN__24[6] __UNCONNECTED_PIN__24[5]
+ __UNCONNECTED_PIN__24[4] __UNCONNECTED_PIN__24[3] __UNCONNECTED_PIN__24[2] __UNCONNECTED_PIN__24[1] __UNCONNECTED_PIN__24[0]
+ __UNCONNECTED_PIN__25[17] __UNCONNECTED_PIN__25[16] __UNCONNECTED_PIN__25[15] __UNCONNECTED_PIN__25[14]
+ __UNCONNECTED_PIN__25[13] __UNCONNECTED_PIN__25[12] __UNCONNECTED_PIN__25[11] __UNCONNECTED_PIN__25[10]
+ __UNCONNECTED_PIN__25[9] __UNCONNECTED_PIN__25[8] __UNCONNECTED_PIN__25[7] __UNCONNECTED_PIN__25[6] __UNCONNECTED_PIN__25[5]
+ __UNCONNECTED_PIN__25[4] __UNCONNECTED_PIN__25[3] __UNCONNECTED_PIN__25[2] __UNCONNECTED_PIN__25[1] __UNCONNECTED_PIN__25[0]
+ __UNCONNECTED_PIN__26[17] __UNCONNECTED_PIN__26[16] __UNCONNECTED_PIN__26[15] __UNCONNECTED_PIN__26[14]
+ __UNCONNECTED_PIN__26[13] __UNCONNECTED_PIN__26[12] __UNCONNECTED_PIN__26[11] __UNCONNECTED_PIN__26[10]
+ __UNCONNECTED_PIN__26[9] __UNCONNECTED_PIN__26[8] __UNCONNECTED_PIN__26[7] __UNCONNECTED_PIN__26[6] __UNCONNECTED_PIN__26[5]
+ __UNCONNECTED_PIN__26[4] __UNCONNECTED_PIN__26[3] __UNCONNECTED_PIN__26[2] __UNCONNECTED_PIN__26[1] __UNCONNECTED_PIN__26[0]
+ __UNCONNECTED_PIN__27[10] __UNCONNECTED_PIN__27[9] __UNCONNECTED_PIN__27[8] __UNCONNECTED_PIN__27[7] __UNCONNECTED_PIN__27[6]
+ __UNCONNECTED_PIN__27[5] __UNCONNECTED_PIN__27[4] __UNCONNECTED_PIN__27[3] __UNCONNECTED_PIN__27[2] __UNCONNECTED_PIN__27[1]
+ __UNCONNECTED_PIN__27[0] __UNCONNECTED_PIN__28[2] __UNCONNECTED_PIN__28[1] __UNCONNECTED_PIN__28[0] __UNCONNECTED_PIN__29[2]
+ __UNCONNECTED_PIN__29[1] __UNCONNECTED_PIN__29[0] __UNCONNECTED_PIN__30 __UNCONNECTED_PIN__31[2] __UNCONNECTED_PIN__31[1]
+ __UNCONNECTED_PIN__31[0] user_analog_project_wrapper
**.ends
