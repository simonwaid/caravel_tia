magic
tech sky130A
magscale 1 2
timestamp 1645630008
<< metal1 >>
rect 886 930 978 966
rect 2144 930 2236 966
rect 3402 930 3494 966
rect 4660 930 4752 966
rect 5918 930 6010 966
rect 7176 930 7268 966
rect 8434 930 8526 966
rect 9692 930 9784 966
rect 10952 932 11040 966
rect 890 680 900 880
rect 980 680 990 880
rect 3390 680 3400 880
rect 3480 680 3490 880
rect 5910 680 5920 880
rect 6000 680 6010 880
rect 8430 680 8440 880
rect 8520 680 8530 880
rect 10950 680 10960 880
rect 11040 680 11050 880
rect -370 110 -360 310
rect -300 110 -290 310
rect 2153 107 2163 307
rect 2223 107 2233 307
rect 4663 107 4673 307
rect 4733 107 4743 307
rect 7183 107 7193 307
rect 7253 107 7263 307
rect 9693 107 9703 307
rect 9763 107 9773 307
rect 12213 107 12223 307
rect 12283 107 12293 307
rect 887 21 977 55
rect 2145 21 2235 55
rect 3403 21 3493 55
rect 4661 21 4751 55
rect 5919 21 6009 55
rect 7177 21 7267 55
rect 8435 21 8525 55
rect 9693 21 9783 55
rect 10951 21 11041 55
<< via1 >>
rect 900 680 980 880
rect 3400 680 3480 880
rect 5920 680 6000 880
rect 8440 680 8520 880
rect 10960 680 11040 880
rect -360 110 -300 310
rect 2163 107 2223 307
rect 4673 107 4733 307
rect 7193 107 7253 307
rect 9703 107 9763 307
rect 12223 107 12283 307
<< metal2 >>
rect 900 880 980 890
rect 3400 880 3480 890
rect 5920 880 6000 890
rect 8440 880 8520 890
rect 10960 880 11040 890
rect -360 680 900 880
rect 980 680 3400 880
rect 3480 680 5920 880
rect 6000 680 8440 880
rect 8520 680 10960 880
rect 11040 680 12280 880
rect 900 670 980 680
rect 3400 670 3480 680
rect 5920 670 6000 680
rect 8440 670 8520 680
rect 10960 670 11040 680
rect -370 310 12290 320
rect -370 110 -360 310
rect -300 307 12290 310
rect -300 110 2163 307
rect -370 107 2163 110
rect 2223 107 4673 307
rect 4733 107 7193 307
rect 7253 107 9703 307
rect 9763 107 12223 307
rect 12283 107 12290 307
rect -370 100 12290 107
rect 2163 97 2223 100
rect 4673 97 4733 100
rect 7193 97 7253 100
rect 9703 97 9763 100
rect 12223 97 12283 100
use sky130_fd_pr__nfet_01v8_HZ8P49  sky130_fd_pr__nfet_01v8_HZ8P49_0
timestamp 1645630008
transform 1 0 5964 0 1 493
box -6457 -610 6457 610
<< end >>
