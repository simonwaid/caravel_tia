* SPICE3 file created from tia_core.ext - technology: sky130A

X0 VN Disable_TIA Disable_TIA_B VN sky130_fd_pr__nfet_01v8 ad=9.6035e+13p pd=6.2292e+08u as=0p ps=0u w=500000u l=1e+06u
X1 VM6D I_Bias1 I_Bias1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.9e+12p ps=4.19e+07u w=2e+06u l=150000u
X2 VM6D I_Bias1 I_Bias1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3 I_Bias1 I_Bias1 VM6D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4 I_Bias1 I_Bias1 VM6D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5 VM6D I_Bias1 I_Bias1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6 VM6D I_Bias1 I_Bias1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7 VM6D I_Bias1 I_Bias1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8 I_Bias1 I_Bias1 VM6D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9 I_Bias1 I_Bias1 VM6D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10 I_Bias1 I_Bias1 VM6D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11 I_Bias1 I_Bias1 VM6D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12 VM6D I_Bias1 I_Bias1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13 VN I_Bias1 VM6D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14 VM6D I_Bias1 VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15 VM6D I_Bias1 VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X16 VN I_Bias1 VM6D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X17 VM6D I_Bias1 VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X18 VN I_Bias1 VM6D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X19 VM5D I_Bias1 Out_1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.412e+13p ps=2.6612e+08u w=2e+06u l=150000u
X20 VM5D I_Bias1 Out_1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X21 Out_1 I_Bias1 VM5D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X22 Out_1 I_Bias1 VM5D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X23 VM5D I_Bias1 Out_1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X24 VM5D I_Bias1 Out_1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X25 VM5D I_Bias1 Out_1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X26 Out_1 I_Bias1 VM5D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X27 Out_1 I_Bias1 VM5D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X28 Out_1 I_Bias1 VM5D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X29 Out_1 I_Bias1 VM5D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X30 VM5D I_Bias1 Out_1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X31 tia_one_tia_0/dis_tran_0/m1_2478_2251# I_Bias1 VM5D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X32 VM5D I_Bias1 tia_one_tia_0/dis_tran_0/m1_2478_2251# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X33 VM5D I_Bias1 tia_one_tia_0/dis_tran_0/m1_2478_2251# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X34 tia_one_tia_0/dis_tran_0/m1_2478_2251# I_Bias1 VM5D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X35 VM5D I_Bias1 tia_one_tia_0/dis_tran_0/m1_2478_2251# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X36 tia_one_tia_0/dis_tran_0/m1_2478_2251# I_Bias1 VM5D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X37 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X38 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X39 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X40 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X41 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X42 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X43 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X44 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X45 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X46 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X47 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X48 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X49 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X50 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X51 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X52 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X53 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X54 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X55 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X56 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X57 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X58 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X59 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X60 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X61 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X62 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X63 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X64 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X65 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X66 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X67 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X68 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X69 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X70 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X71 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X72 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X73 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X74 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X75 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X76 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X77 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X78 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X79 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X80 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X81 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X82 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X83 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X84 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X85 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X86 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X87 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X88 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X89 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X90 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X91 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X92 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X93 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X94 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X95 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X96 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X97 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X98 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X99 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X100 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X101 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X102 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X103 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X104 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X105 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X106 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X107 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X108 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X109 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X110 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X111 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X112 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X113 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X114 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X115 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X116 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X117 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X118 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X119 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X120 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X121 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X122 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X123 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X124 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X125 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X126 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X127 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X128 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X129 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X130 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X131 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X132 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X133 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X134 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X135 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X136 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X137 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=4.3065e+13p pd=3.405e+08u as=1.856e+13p ps=1.4656e+08u w=2e+06u l=200000u
X138 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X139 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X140 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X141 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X142 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X143 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X144 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X145 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X146 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X147 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X148 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X149 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X150 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X151 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X152 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X153 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X154 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X155 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X156 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X157 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X158 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X159 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X160 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X161 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X162 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X163 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X164 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X165 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X166 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X167 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X168 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X169 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X170 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X171 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X172 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X173 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X174 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X175 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X176 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X177 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X178 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X179 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X180 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X181 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X182 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X183 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X184 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X185 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X186 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X187 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X188 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X189 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X190 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X191 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X192 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X193 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X194 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X195 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X196 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X197 VPP tia_one_tia_0/sky130_fd_pr__cap_mim_m3_2_ZWVPUJ_0/m4_n2851_n1900# sky130_fd_pr__cap_mim_m3_2 l=1.8e+07u w=2.5e+07u
X198 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X199 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X200 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X201 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X202 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X203 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X204 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X205 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X206 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X207 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X208 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X209 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X210 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X211 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X212 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X213 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X214 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X215 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X216 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X217 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X218 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X219 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X220 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X221 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X222 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X223 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X224 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X225 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X226 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X227 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X228 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X229 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X230 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X231 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X232 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X233 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X234 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X235 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X236 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X237 tia_one_tia_0/dis_tran_0/m1_2478_2251# Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X238 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X239 tia_one_tia_0/dis_tran_0/m1_2478_2251# Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X240 VM28D Disable_TIA_B tia_one_tia_0/dis_tran_0/m1_2478_2251# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X241 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X242 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X243 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X244 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X245 tia_one_tia_0/dis_tran_0/m1_2478_2251# Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X246 VM28D Disable_TIA_B tia_one_tia_0/dis_tran_0/m1_2478_2251# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X247 tia_one_tia_0/dis_tran_0/m1_2478_2251# Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X248 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X249 VM28D Disable_TIA_B tia_one_tia_0/dis_tran_0/m1_2478_2251# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X250 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X251 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X252 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X253 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X254 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X255 VM28D Disable_TIA_B tia_one_tia_0/dis_tran_0/m1_2478_2251# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X256 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X257 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X258 tia_one_tia_0/dis_tran_0/m1_2478_2251# Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X259 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X260 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X261 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X262 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X263 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X264 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X265 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X266 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X267 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X268 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X269 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X270 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X271 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X272 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X273 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X274 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X275 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X276 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X277 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X278 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X279 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X280 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X281 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X282 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X283 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X284 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X285 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X286 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X287 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X288 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X289 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X290 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X291 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X292 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X293 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X294 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X295 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X296 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X297 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X298 Out_2 VN VPP VPP sky130_fd_pr__pfet_01v8 ad=3.48e+12p pd=2.748e+07u as=0p ps=0u w=2e+06u l=500000u
X299 Out_2 VN VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X300 VPP VN Out_2 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X301 VPP VN Out_2 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X302 Out_2 VN VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X303 Out_2 VN VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X304 Out_2 VN VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X305 VPP VN Out_2 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X306 VPP VN Out_2 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X307 VPP VN Out_2 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X308 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=3.56368e+13p pd=5.4965e+07u as=9.28e+12p ps=7.328e+07u w=2e+06u l=200000u
X309 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X310 Out_2 Out_1 Input Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X311 Out_2 Out_1 Input Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X312 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X313 Out_2 Out_1 Input Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X314 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X315 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X316 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X317 Out_2 Out_1 Input Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X318 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X319 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X320 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X321 Out_2 Out_1 Input Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X322 Out_2 Out_1 Input Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X323 Out_2 Out_1 Input Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X324 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X325 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X326 Out_2 Out_1 Input Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X327 Out_2 Out_1 Input Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X328 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X329 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X330 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X331 Out_2 Out_1 Input Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X332 Out_2 Out_1 Input Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X333 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X334 Out_2 Out_1 Input Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X335 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X336 Out_2 Out_1 Input Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X337 Out_2 Out_1 Input Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X338 tia_one_tia_1/tia_cur_mirror_0/m1_71_130# I_Bias1 tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X339 tia_one_tia_1/tia_cur_mirror_0/m1_71_130# I_Bias1 tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X340 tia_one_tia_1/m1_1540_1550# I_Bias1 tia_one_tia_1/tia_cur_mirror_0/m1_71_130# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X341 tia_one_tia_1/m1_1540_1550# I_Bias1 tia_one_tia_1/tia_cur_mirror_0/m1_71_130# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X342 tia_one_tia_1/tia_cur_mirror_0/m1_71_130# I_Bias1 tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X343 tia_one_tia_1/tia_cur_mirror_0/m1_71_130# I_Bias1 tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X344 tia_one_tia_1/tia_cur_mirror_0/m1_71_130# I_Bias1 tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X345 tia_one_tia_1/m1_1540_1550# I_Bias1 tia_one_tia_1/tia_cur_mirror_0/m1_71_130# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X346 tia_one_tia_1/m1_1540_1550# I_Bias1 tia_one_tia_1/tia_cur_mirror_0/m1_71_130# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X347 tia_one_tia_1/m1_1540_1550# I_Bias1 tia_one_tia_1/tia_cur_mirror_0/m1_71_130# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X348 tia_one_tia_1/m1_1540_1550# I_Bias1 tia_one_tia_1/tia_cur_mirror_0/m1_71_130# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X349 tia_one_tia_1/tia_cur_mirror_0/m1_71_130# I_Bias1 tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X350 VN I_Bias1 tia_one_tia_1/tia_cur_mirror_0/m1_71_130# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X351 tia_one_tia_1/tia_cur_mirror_0/m1_71_130# I_Bias1 VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X352 tia_one_tia_1/tia_cur_mirror_0/m1_71_130# I_Bias1 VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X353 VN I_Bias1 tia_one_tia_1/tia_cur_mirror_0/m1_71_130# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X354 tia_one_tia_1/tia_cur_mirror_0/m1_71_130# I_Bias1 VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X355 VN I_Bias1 tia_one_tia_1/tia_cur_mirror_0/m1_71_130# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X356 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X357 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X358 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X359 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X360 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X361 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X362 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X363 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X364 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X365 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X366 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X367 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X368 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X369 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X370 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X371 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X372 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X373 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X374 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X375 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X376 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X377 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X378 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X379 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X380 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X381 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X382 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X383 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X384 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X385 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X386 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X387 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X388 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X389 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X390 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X391 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X392 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X393 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X394 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X395 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X396 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X397 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X398 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X399 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X400 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X401 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X402 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X403 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X404 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X405 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X406 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X407 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X408 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X409 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X410 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X411 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X412 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X413 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X414 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X415 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X416 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X417 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X418 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X419 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X420 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X421 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X422 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X423 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X424 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X425 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X426 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X427 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X428 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X429 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X430 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X431 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X432 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X433 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X434 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X435 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X436 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X437 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X438 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X439 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X440 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X441 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X442 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X443 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X444 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X445 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X446 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X447 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X448 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X449 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X450 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X451 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X452 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X453 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X454 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X455 VM40D w_2300_n7574# tia_one_tia_1/m1_1540_1550# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X456 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X457 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X458 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X459 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X460 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X461 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X462 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X463 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X464 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X465 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X466 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X467 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X468 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X469 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X470 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X471 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X472 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X473 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X474 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X475 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X476 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X477 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X478 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X479 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X480 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X481 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X482 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X483 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X484 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X485 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X486 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X487 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X488 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X489 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X490 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X491 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X492 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X493 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X494 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X495 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X496 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X497 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X498 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X499 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X500 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X501 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X502 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X503 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X504 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X505 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X506 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X507 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X508 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X509 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X510 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X511 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X512 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X513 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X514 tia_one_tia_1/m1_1540_1550# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X515 VPP w_2300_n7574# tia_one_tia_1/m1_1540_1550# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X516 VPP tia_one_tia_1/sky130_fd_pr__cap_mim_m3_2_ZWVPUJ_0/m4_n2851_n1900# sky130_fd_pr__cap_mim_m3_2 l=1.8e+07u w=2.5e+07u
X517 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X518 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X519 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X520 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X521 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X522 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X523 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X524 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X525 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X526 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X527 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X528 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X529 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X530 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X531 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X532 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X533 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X534 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X535 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X536 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X537 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X538 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X539 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X540 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X541 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X542 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X543 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X544 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X545 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X546 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X547 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X548 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X549 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X550 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X551 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X552 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X553 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X554 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X555 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X556 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X557 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X558 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X559 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X560 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X561 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X562 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X563 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X564 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X565 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X566 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X567 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X568 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X569 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X570 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X571 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X572 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X573 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X574 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X575 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X576 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X577 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X578 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X579 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X580 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X581 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X582 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X583 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X584 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X585 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X586 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X587 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X588 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X589 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X590 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X591 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X592 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X593 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X594 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X595 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X596 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X597 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X598 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X599 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X600 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X601 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X602 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X603 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X604 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X605 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X606 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X607 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X608 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X609 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X610 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X611 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X612 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X613 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X614 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X615 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X616 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X617 m3_2920_n6050# VN VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X618 m3_2920_n6050# VN VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X619 VPP VN m3_2920_n6050# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X620 VPP VN m3_2920_n6050# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X621 m3_2920_n6050# VN VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X622 m3_2920_n6050# VN VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X623 m3_2920_n6050# VN VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X624 VPP VN m3_2920_n6050# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X625 VPP VN m3_2920_n6050# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X626 VPP VN m3_2920_n6050# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X627 w_2300_n7574# tia_one_tia_1/m1_1540_1550# m3_2920_n6050# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X628 w_2300_n7574# tia_one_tia_1/m1_1540_1550# m3_2920_n6050# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X629 m3_2920_n6050# tia_one_tia_1/m1_1540_1550# w_2300_n7574# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X630 m3_2920_n6050# tia_one_tia_1/m1_1540_1550# w_2300_n7574# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X631 w_2300_n7574# tia_one_tia_1/m1_1540_1550# m3_2920_n6050# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X632 m3_2920_n6050# tia_one_tia_1/m1_1540_1550# w_2300_n7574# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X633 w_2300_n7574# tia_one_tia_1/m1_1540_1550# m3_2920_n6050# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X634 w_2300_n7574# tia_one_tia_1/m1_1540_1550# m3_2920_n6050# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X635 w_2300_n7574# tia_one_tia_1/m1_1540_1550# m3_2920_n6050# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X636 m3_2920_n6050# tia_one_tia_1/m1_1540_1550# w_2300_n7574# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X637 w_2300_n7574# tia_one_tia_1/m1_1540_1550# m3_2920_n6050# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X638 w_2300_n7574# tia_one_tia_1/m1_1540_1550# m3_2920_n6050# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X639 w_2300_n7574# tia_one_tia_1/m1_1540_1550# m3_2920_n6050# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X640 m3_2920_n6050# tia_one_tia_1/m1_1540_1550# w_2300_n7574# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X641 m3_2920_n6050# tia_one_tia_1/m1_1540_1550# w_2300_n7574# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X642 m3_2920_n6050# tia_one_tia_1/m1_1540_1550# w_2300_n7574# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X643 w_2300_n7574# tia_one_tia_1/m1_1540_1550# m3_2920_n6050# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X644 w_2300_n7574# tia_one_tia_1/m1_1540_1550# m3_2920_n6050# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X645 m3_2920_n6050# tia_one_tia_1/m1_1540_1550# w_2300_n7574# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X646 m3_2920_n6050# tia_one_tia_1/m1_1540_1550# w_2300_n7574# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X647 w_2300_n7574# tia_one_tia_1/m1_1540_1550# m3_2920_n6050# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X648 w_2300_n7574# tia_one_tia_1/m1_1540_1550# m3_2920_n6050# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X649 w_2300_n7574# tia_one_tia_1/m1_1540_1550# m3_2920_n6050# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X650 m3_2920_n6050# tia_one_tia_1/m1_1540_1550# w_2300_n7574# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X651 m3_2920_n6050# tia_one_tia_1/m1_1540_1550# w_2300_n7574# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X652 w_2300_n7574# tia_one_tia_1/m1_1540_1550# m3_2920_n6050# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X653 m3_2920_n6050# tia_one_tia_1/m1_1540_1550# w_2300_n7574# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X654 w_2300_n7574# tia_one_tia_1/m1_1540_1550# m3_2920_n6050# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X655 m3_2920_n6050# tia_one_tia_1/m1_1540_1550# w_2300_n7574# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X656 m3_2920_n6050# tia_one_tia_1/m1_1540_1550# w_2300_n7574# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X657 VPP Disable_TIA Disable_TIA_B VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=1e+06u
X658 VN I_Bias1 sky130_fd_pr__cap_mim_m3_1 l=1.2e+07u w=1.5e+07u
X659 VN I_Bias1 sky130_fd_pr__cap_mim_m3_1 l=1.2e+07u w=1.5e+07u
X660 Disable_TIA_B VN VN sky130_fd_pr__cap_var_lvt pd=0u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X661 Disable_TIA_B VN VN sky130_fd_pr__cap_var_lvt pd=0u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X662 Disable_TIA_B VN VN sky130_fd_pr__cap_var_lvt pd=0u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X663 Disable_TIA_B VN VN sky130_fd_pr__cap_var_lvt pd=0u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X664 Disable_TIA_B VN VN sky130_fd_pr__cap_var_lvt pd=0u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X665 VPP VN sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X666 VPP VN sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X667 I_Bias1 Disable_TIA VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X668 VN Disable_TIA I_Bias1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X669 VN Disable_TIA I_Bias1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X670 VN Disable_TIA I_Bias1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X671 I_Bias1 Disable_TIA VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
