magic
tech sky130A
magscale 1 2
timestamp 1646921651
<< nwell >>
rect -683 -1373 683 1373
<< pmos >>
rect -487 754 -287 1154
rect -229 754 -29 1154
rect 29 754 229 1154
rect 287 754 487 1154
rect -487 118 -287 518
rect -229 118 -29 518
rect 29 118 229 518
rect 287 118 487 518
rect -487 -518 -287 -118
rect -229 -518 -29 -118
rect 29 -518 229 -118
rect 287 -518 487 -118
rect -487 -1154 -287 -754
rect -229 -1154 -29 -754
rect 29 -1154 229 -754
rect 287 -1154 487 -754
<< pdiff >>
rect -545 1142 -487 1154
rect -545 766 -533 1142
rect -499 766 -487 1142
rect -545 754 -487 766
rect -287 1142 -229 1154
rect -287 766 -275 1142
rect -241 766 -229 1142
rect -287 754 -229 766
rect -29 1142 29 1154
rect -29 766 -17 1142
rect 17 766 29 1142
rect -29 754 29 766
rect 229 1142 287 1154
rect 229 766 241 1142
rect 275 766 287 1142
rect 229 754 287 766
rect 487 1142 545 1154
rect 487 766 499 1142
rect 533 766 545 1142
rect 487 754 545 766
rect -545 506 -487 518
rect -545 130 -533 506
rect -499 130 -487 506
rect -545 118 -487 130
rect -287 506 -229 518
rect -287 130 -275 506
rect -241 130 -229 506
rect -287 118 -229 130
rect -29 506 29 518
rect -29 130 -17 506
rect 17 130 29 506
rect -29 118 29 130
rect 229 506 287 518
rect 229 130 241 506
rect 275 130 287 506
rect 229 118 287 130
rect 487 506 545 518
rect 487 130 499 506
rect 533 130 545 506
rect 487 118 545 130
rect -545 -130 -487 -118
rect -545 -506 -533 -130
rect -499 -506 -487 -130
rect -545 -518 -487 -506
rect -287 -130 -229 -118
rect -287 -506 -275 -130
rect -241 -506 -229 -130
rect -287 -518 -229 -506
rect -29 -130 29 -118
rect -29 -506 -17 -130
rect 17 -506 29 -130
rect -29 -518 29 -506
rect 229 -130 287 -118
rect 229 -506 241 -130
rect 275 -506 287 -130
rect 229 -518 287 -506
rect 487 -130 545 -118
rect 487 -506 499 -130
rect 533 -506 545 -130
rect 487 -518 545 -506
rect -545 -766 -487 -754
rect -545 -1142 -533 -766
rect -499 -1142 -487 -766
rect -545 -1154 -487 -1142
rect -287 -766 -229 -754
rect -287 -1142 -275 -766
rect -241 -1142 -229 -766
rect -287 -1154 -229 -1142
rect -29 -766 29 -754
rect -29 -1142 -17 -766
rect 17 -1142 29 -766
rect -29 -1154 29 -1142
rect 229 -766 287 -754
rect 229 -1142 241 -766
rect 275 -1142 287 -766
rect 229 -1154 287 -1142
rect 487 -766 545 -754
rect 487 -1142 499 -766
rect 533 -1142 545 -766
rect 487 -1154 545 -1142
<< pdiffc >>
rect -533 766 -499 1142
rect -275 766 -241 1142
rect -17 766 17 1142
rect 241 766 275 1142
rect 499 766 533 1142
rect -533 130 -499 506
rect -275 130 -241 506
rect -17 130 17 506
rect 241 130 275 506
rect 499 130 533 506
rect -533 -506 -499 -130
rect -275 -506 -241 -130
rect -17 -506 17 -130
rect 241 -506 275 -130
rect 499 -506 533 -130
rect -533 -1142 -499 -766
rect -275 -1142 -241 -766
rect -17 -1142 17 -766
rect 241 -1142 275 -766
rect 499 -1142 533 -766
<< nsubdiff >>
rect -647 1303 -551 1337
rect 551 1303 647 1337
rect -647 1241 -613 1303
rect 613 1241 647 1303
rect -647 -1303 -613 -1241
rect 613 -1303 647 -1241
rect -647 -1337 -551 -1303
rect 551 -1337 647 -1303
<< nsubdiffcont >>
rect -551 1303 551 1337
rect -647 -1241 -613 1241
rect 613 -1241 647 1241
rect -551 -1337 551 -1303
<< poly >>
rect -487 1235 -287 1251
rect -487 1201 -471 1235
rect -303 1201 -287 1235
rect -487 1154 -287 1201
rect -229 1235 -29 1251
rect -229 1201 -213 1235
rect -45 1201 -29 1235
rect -229 1154 -29 1201
rect 29 1235 229 1251
rect 29 1201 45 1235
rect 213 1201 229 1235
rect 29 1154 229 1201
rect 287 1235 487 1251
rect 287 1201 303 1235
rect 471 1201 487 1235
rect 287 1154 487 1201
rect -487 707 -287 754
rect -487 673 -471 707
rect -303 673 -287 707
rect -487 657 -287 673
rect -229 707 -29 754
rect -229 673 -213 707
rect -45 673 -29 707
rect -229 657 -29 673
rect 29 707 229 754
rect 29 673 45 707
rect 213 673 229 707
rect 29 657 229 673
rect 287 707 487 754
rect 287 673 303 707
rect 471 673 487 707
rect 287 657 487 673
rect -487 599 -287 615
rect -487 565 -471 599
rect -303 565 -287 599
rect -487 518 -287 565
rect -229 599 -29 615
rect -229 565 -213 599
rect -45 565 -29 599
rect -229 518 -29 565
rect 29 599 229 615
rect 29 565 45 599
rect 213 565 229 599
rect 29 518 229 565
rect 287 599 487 615
rect 287 565 303 599
rect 471 565 487 599
rect 287 518 487 565
rect -487 71 -287 118
rect -487 37 -471 71
rect -303 37 -287 71
rect -487 21 -287 37
rect -229 71 -29 118
rect -229 37 -213 71
rect -45 37 -29 71
rect -229 21 -29 37
rect 29 71 229 118
rect 29 37 45 71
rect 213 37 229 71
rect 29 21 229 37
rect 287 71 487 118
rect 287 37 303 71
rect 471 37 487 71
rect 287 21 487 37
rect -487 -37 -287 -21
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -487 -118 -287 -71
rect -229 -37 -29 -21
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect -229 -118 -29 -71
rect 29 -37 229 -21
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 29 -118 229 -71
rect 287 -37 487 -21
rect 287 -71 303 -37
rect 471 -71 487 -37
rect 287 -118 487 -71
rect -487 -565 -287 -518
rect -487 -599 -471 -565
rect -303 -599 -287 -565
rect -487 -615 -287 -599
rect -229 -565 -29 -518
rect -229 -599 -213 -565
rect -45 -599 -29 -565
rect -229 -615 -29 -599
rect 29 -565 229 -518
rect 29 -599 45 -565
rect 213 -599 229 -565
rect 29 -615 229 -599
rect 287 -565 487 -518
rect 287 -599 303 -565
rect 471 -599 487 -565
rect 287 -615 487 -599
rect -487 -673 -287 -657
rect -487 -707 -471 -673
rect -303 -707 -287 -673
rect -487 -754 -287 -707
rect -229 -673 -29 -657
rect -229 -707 -213 -673
rect -45 -707 -29 -673
rect -229 -754 -29 -707
rect 29 -673 229 -657
rect 29 -707 45 -673
rect 213 -707 229 -673
rect 29 -754 229 -707
rect 287 -673 487 -657
rect 287 -707 303 -673
rect 471 -707 487 -673
rect 287 -754 487 -707
rect -487 -1201 -287 -1154
rect -487 -1235 -471 -1201
rect -303 -1235 -287 -1201
rect -487 -1251 -287 -1235
rect -229 -1201 -29 -1154
rect -229 -1235 -213 -1201
rect -45 -1235 -29 -1201
rect -229 -1251 -29 -1235
rect 29 -1201 229 -1154
rect 29 -1235 45 -1201
rect 213 -1235 229 -1201
rect 29 -1251 229 -1235
rect 287 -1201 487 -1154
rect 287 -1235 303 -1201
rect 471 -1235 487 -1201
rect 287 -1251 487 -1235
<< polycont >>
rect -471 1201 -303 1235
rect -213 1201 -45 1235
rect 45 1201 213 1235
rect 303 1201 471 1235
rect -471 673 -303 707
rect -213 673 -45 707
rect 45 673 213 707
rect 303 673 471 707
rect -471 565 -303 599
rect -213 565 -45 599
rect 45 565 213 599
rect 303 565 471 599
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect -471 -599 -303 -565
rect -213 -599 -45 -565
rect 45 -599 213 -565
rect 303 -599 471 -565
rect -471 -707 -303 -673
rect -213 -707 -45 -673
rect 45 -707 213 -673
rect 303 -707 471 -673
rect -471 -1235 -303 -1201
rect -213 -1235 -45 -1201
rect 45 -1235 213 -1201
rect 303 -1235 471 -1201
<< locali >>
rect -647 1303 -551 1337
rect 551 1303 647 1337
rect -647 1241 -613 1303
rect 613 1241 647 1303
rect -487 1201 -471 1235
rect -303 1201 -287 1235
rect -229 1201 -213 1235
rect -45 1201 -29 1235
rect 29 1201 45 1235
rect 213 1201 229 1235
rect 287 1201 303 1235
rect 471 1201 487 1235
rect -533 1142 -499 1158
rect -533 750 -499 766
rect -275 1142 -241 1158
rect -275 750 -241 766
rect -17 1142 17 1158
rect -17 750 17 766
rect 241 1142 275 1158
rect 241 750 275 766
rect 499 1142 533 1158
rect 499 750 533 766
rect -487 673 -471 707
rect -303 673 -287 707
rect -229 673 -213 707
rect -45 673 -29 707
rect 29 673 45 707
rect 213 673 229 707
rect 287 673 303 707
rect 471 673 487 707
rect -487 565 -471 599
rect -303 565 -287 599
rect -229 565 -213 599
rect -45 565 -29 599
rect 29 565 45 599
rect 213 565 229 599
rect 287 565 303 599
rect 471 565 487 599
rect -533 506 -499 522
rect -533 114 -499 130
rect -275 506 -241 522
rect -275 114 -241 130
rect -17 506 17 522
rect -17 114 17 130
rect 241 506 275 522
rect 241 114 275 130
rect 499 506 533 522
rect 499 114 533 130
rect -487 37 -471 71
rect -303 37 -287 71
rect -229 37 -213 71
rect -45 37 -29 71
rect 29 37 45 71
rect 213 37 229 71
rect 287 37 303 71
rect 471 37 487 71
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 287 -71 303 -37
rect 471 -71 487 -37
rect -533 -130 -499 -114
rect -533 -522 -499 -506
rect -275 -130 -241 -114
rect -275 -522 -241 -506
rect -17 -130 17 -114
rect -17 -522 17 -506
rect 241 -130 275 -114
rect 241 -522 275 -506
rect 499 -130 533 -114
rect 499 -522 533 -506
rect -487 -599 -471 -565
rect -303 -599 -287 -565
rect -229 -599 -213 -565
rect -45 -599 -29 -565
rect 29 -599 45 -565
rect 213 -599 229 -565
rect 287 -599 303 -565
rect 471 -599 487 -565
rect -487 -707 -471 -673
rect -303 -707 -287 -673
rect -229 -707 -213 -673
rect -45 -707 -29 -673
rect 29 -707 45 -673
rect 213 -707 229 -673
rect 287 -707 303 -673
rect 471 -707 487 -673
rect -533 -766 -499 -750
rect -533 -1158 -499 -1142
rect -275 -766 -241 -750
rect -275 -1158 -241 -1142
rect -17 -766 17 -750
rect -17 -1158 17 -1142
rect 241 -766 275 -750
rect 241 -1158 275 -1142
rect 499 -766 533 -750
rect 499 -1158 533 -1142
rect -487 -1235 -471 -1201
rect -303 -1235 -287 -1201
rect -229 -1235 -213 -1201
rect -45 -1235 -29 -1201
rect 29 -1235 45 -1201
rect 213 -1235 229 -1201
rect 287 -1235 303 -1201
rect 471 -1235 487 -1201
rect -647 -1303 -613 -1241
rect 613 -1303 647 -1241
rect -647 -1337 -551 -1303
rect 551 -1337 647 -1303
<< viali >>
rect -471 1201 -303 1235
rect -213 1201 -45 1235
rect 45 1201 213 1235
rect 303 1201 471 1235
rect -533 766 -499 1142
rect -275 766 -241 1142
rect -17 766 17 1142
rect 241 766 275 1142
rect 499 766 533 1142
rect -471 673 -303 707
rect -213 673 -45 707
rect 45 673 213 707
rect 303 673 471 707
rect -471 565 -303 599
rect -213 565 -45 599
rect 45 565 213 599
rect 303 565 471 599
rect -533 130 -499 506
rect -275 130 -241 506
rect -17 130 17 506
rect 241 130 275 506
rect 499 130 533 506
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect -533 -506 -499 -130
rect -275 -506 -241 -130
rect -17 -506 17 -130
rect 241 -506 275 -130
rect 499 -506 533 -130
rect -471 -599 -303 -565
rect -213 -599 -45 -565
rect 45 -599 213 -565
rect 303 -599 471 -565
rect -471 -707 -303 -673
rect -213 -707 -45 -673
rect 45 -707 213 -673
rect 303 -707 471 -673
rect -533 -1142 -499 -766
rect -275 -1142 -241 -766
rect -17 -1142 17 -766
rect 241 -1142 275 -766
rect 499 -1142 533 -766
rect -471 -1235 -303 -1201
rect -213 -1235 -45 -1201
rect 45 -1235 213 -1201
rect 303 -1235 471 -1201
<< metal1 >>
rect -483 1235 -291 1241
rect -483 1201 -471 1235
rect -303 1201 -291 1235
rect -483 1195 -291 1201
rect -225 1235 -33 1241
rect -225 1201 -213 1235
rect -45 1201 -33 1235
rect -225 1195 -33 1201
rect 33 1235 225 1241
rect 33 1201 45 1235
rect 213 1201 225 1235
rect 33 1195 225 1201
rect 291 1235 483 1241
rect 291 1201 303 1235
rect 471 1201 483 1235
rect 291 1195 483 1201
rect -539 1142 -493 1154
rect -539 766 -533 1142
rect -499 766 -493 1142
rect -539 754 -493 766
rect -281 1142 -235 1154
rect -281 766 -275 1142
rect -241 766 -235 1142
rect -281 754 -235 766
rect -23 1142 23 1154
rect -23 766 -17 1142
rect 17 766 23 1142
rect -23 754 23 766
rect 235 1142 281 1154
rect 235 766 241 1142
rect 275 766 281 1142
rect 235 754 281 766
rect 493 1142 539 1154
rect 493 766 499 1142
rect 533 766 539 1142
rect 493 754 539 766
rect -483 707 -291 713
rect -483 673 -471 707
rect -303 673 -291 707
rect -483 667 -291 673
rect -225 707 -33 713
rect -225 673 -213 707
rect -45 673 -33 707
rect -225 667 -33 673
rect 33 707 225 713
rect 33 673 45 707
rect 213 673 225 707
rect 33 667 225 673
rect 291 707 483 713
rect 291 673 303 707
rect 471 673 483 707
rect 291 667 483 673
rect -483 599 -291 605
rect -483 565 -471 599
rect -303 565 -291 599
rect -483 559 -291 565
rect -225 599 -33 605
rect -225 565 -213 599
rect -45 565 -33 599
rect -225 559 -33 565
rect 33 599 225 605
rect 33 565 45 599
rect 213 565 225 599
rect 33 559 225 565
rect 291 599 483 605
rect 291 565 303 599
rect 471 565 483 599
rect 291 559 483 565
rect -539 506 -493 518
rect -539 130 -533 506
rect -499 130 -493 506
rect -539 118 -493 130
rect -281 506 -235 518
rect -281 130 -275 506
rect -241 130 -235 506
rect -281 118 -235 130
rect -23 506 23 518
rect -23 130 -17 506
rect 17 130 23 506
rect -23 118 23 130
rect 235 506 281 518
rect 235 130 241 506
rect 275 130 281 506
rect 235 118 281 130
rect 493 506 539 518
rect 493 130 499 506
rect 533 130 539 506
rect 493 118 539 130
rect -483 71 -291 77
rect -483 37 -471 71
rect -303 37 -291 71
rect -483 31 -291 37
rect -225 71 -33 77
rect -225 37 -213 71
rect -45 37 -33 71
rect -225 31 -33 37
rect 33 71 225 77
rect 33 37 45 71
rect 213 37 225 71
rect 33 31 225 37
rect 291 71 483 77
rect 291 37 303 71
rect 471 37 483 71
rect 291 31 483 37
rect -483 -37 -291 -31
rect -483 -71 -471 -37
rect -303 -71 -291 -37
rect -483 -77 -291 -71
rect -225 -37 -33 -31
rect -225 -71 -213 -37
rect -45 -71 -33 -37
rect -225 -77 -33 -71
rect 33 -37 225 -31
rect 33 -71 45 -37
rect 213 -71 225 -37
rect 33 -77 225 -71
rect 291 -37 483 -31
rect 291 -71 303 -37
rect 471 -71 483 -37
rect 291 -77 483 -71
rect -539 -130 -493 -118
rect -539 -506 -533 -130
rect -499 -506 -493 -130
rect -539 -518 -493 -506
rect -281 -130 -235 -118
rect -281 -506 -275 -130
rect -241 -506 -235 -130
rect -281 -518 -235 -506
rect -23 -130 23 -118
rect -23 -506 -17 -130
rect 17 -506 23 -130
rect -23 -518 23 -506
rect 235 -130 281 -118
rect 235 -506 241 -130
rect 275 -506 281 -130
rect 235 -518 281 -506
rect 493 -130 539 -118
rect 493 -506 499 -130
rect 533 -506 539 -130
rect 493 -518 539 -506
rect -483 -565 -291 -559
rect -483 -599 -471 -565
rect -303 -599 -291 -565
rect -483 -605 -291 -599
rect -225 -565 -33 -559
rect -225 -599 -213 -565
rect -45 -599 -33 -565
rect -225 -605 -33 -599
rect 33 -565 225 -559
rect 33 -599 45 -565
rect 213 -599 225 -565
rect 33 -605 225 -599
rect 291 -565 483 -559
rect 291 -599 303 -565
rect 471 -599 483 -565
rect 291 -605 483 -599
rect -483 -673 -291 -667
rect -483 -707 -471 -673
rect -303 -707 -291 -673
rect -483 -713 -291 -707
rect -225 -673 -33 -667
rect -225 -707 -213 -673
rect -45 -707 -33 -673
rect -225 -713 -33 -707
rect 33 -673 225 -667
rect 33 -707 45 -673
rect 213 -707 225 -673
rect 33 -713 225 -707
rect 291 -673 483 -667
rect 291 -707 303 -673
rect 471 -707 483 -673
rect 291 -713 483 -707
rect -539 -766 -493 -754
rect -539 -1142 -533 -766
rect -499 -1142 -493 -766
rect -539 -1154 -493 -1142
rect -281 -766 -235 -754
rect -281 -1142 -275 -766
rect -241 -1142 -235 -766
rect -281 -1154 -235 -1142
rect -23 -766 23 -754
rect -23 -1142 -17 -766
rect 17 -1142 23 -766
rect -23 -1154 23 -1142
rect 235 -766 281 -754
rect 235 -1142 241 -766
rect 275 -1142 281 -766
rect 235 -1154 281 -1142
rect 493 -766 539 -754
rect 493 -1142 499 -766
rect 533 -1142 539 -766
rect 493 -1154 539 -1142
rect -483 -1201 -291 -1195
rect -483 -1235 -471 -1201
rect -303 -1235 -291 -1201
rect -483 -1241 -291 -1235
rect -225 -1201 -33 -1195
rect -225 -1235 -213 -1201
rect -45 -1235 -33 -1201
rect -225 -1241 -33 -1235
rect 33 -1201 225 -1195
rect 33 -1235 45 -1201
rect 213 -1235 225 -1201
rect 33 -1241 225 -1235
rect 291 -1201 483 -1195
rect 291 -1235 303 -1201
rect 471 -1235 483 -1201
rect 291 -1241 483 -1235
<< properties >>
string FIXED_BBOX -630 -1320 630 1320
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 1 m 4 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
