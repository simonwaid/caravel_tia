magic
tech sky130A
timestamp 1646921651
<< pwell >>
rect -148 -130 148 130
<< nmos >>
rect -50 -25 50 25
<< ndiff >>
rect -79 19 -50 25
rect -79 -19 -73 19
rect -56 -19 -50 19
rect -79 -25 -50 -19
rect 50 19 79 25
rect 50 -19 56 19
rect 73 -19 79 19
rect 50 -25 79 -19
<< ndiffc >>
rect -73 -19 -56 19
rect 56 -19 73 19
<< psubdiff >>
rect -130 95 -82 112
rect 82 95 130 112
rect -130 64 -113 95
rect 113 64 130 95
rect -130 -95 -113 -64
rect 113 -95 130 -64
rect -130 -112 -82 -95
rect 82 -112 130 -95
<< psubdiffcont >>
rect -82 95 82 112
rect -130 -64 -113 64
rect 113 -64 130 64
rect -82 -112 82 -95
<< poly >>
rect -50 61 50 69
rect -50 44 -42 61
rect 42 44 50 61
rect -50 25 50 44
rect -50 -44 50 -25
rect -50 -61 -42 -44
rect 42 -61 50 -44
rect -50 -69 50 -61
<< polycont >>
rect -42 44 42 61
rect -42 -61 42 -44
<< locali >>
rect -130 95 -82 112
rect 82 95 130 112
rect -130 64 -113 95
rect 113 64 130 95
rect -50 44 -42 61
rect 42 44 50 61
rect -73 19 -56 27
rect -73 -27 -56 -19
rect 56 19 73 27
rect 56 -27 73 -19
rect -50 -61 -42 -44
rect 42 -61 50 -44
rect -130 -95 -113 -64
rect 113 -95 130 -64
rect -130 -112 -82 -95
rect 82 -112 130 -95
<< viali >>
rect -42 44 42 61
rect -73 -19 -56 19
rect 56 -19 73 19
rect -42 -61 42 -44
<< metal1 >>
rect -48 61 48 64
rect -48 44 -42 61
rect 42 44 48 61
rect -48 41 48 44
rect -76 19 -53 25
rect -76 -19 -73 19
rect -56 -19 -53 19
rect -76 -25 -53 -19
rect 53 19 76 25
rect 53 -19 56 19
rect 73 -19 76 19
rect 53 -25 76 -19
rect -48 -44 48 -41
rect -48 -61 -42 -44
rect 42 -61 48 -44
rect -48 -64 48 -61
<< properties >>
string FIXED_BBOX -121 -103 121 103
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 1 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
