magic
tech sky130A
magscale 1 2
timestamp 1647269090
<< locali >>
rect 3230 -2570 5340 -2130
rect 4108 -7934 4420 -7920
rect 3740 -7940 4420 -7934
rect 3300 -9460 3420 -8660
rect 4800 -8730 5340 -2570
rect 4800 -8740 5390 -8730
rect 4800 -8750 5370 -8740
rect 3300 -9470 4420 -9460
rect 5200 -9470 5370 -8750
rect 5960 -9310 6070 -9150
rect 5970 -9320 6070 -9310
rect 5980 -9470 6070 -9320
rect 1340 -9740 6090 -9470
rect 1340 -9750 4800 -9740
rect 1340 -11100 1510 -9750
rect 2160 -11100 2540 -9750
rect 3070 -11100 3450 -9750
rect 4000 -11100 4380 -9750
rect 4910 -11100 5310 -9740
rect 5840 -11090 5960 -9750
rect 6620 -10320 6670 -10200
rect 5970 -11040 6240 -10600
rect 6610 -10880 6710 -10760
rect 1340 -11280 5970 -11100
<< viali >>
rect 6670 -10320 6760 -10200
<< metal1 >>
rect 4100 1996 4660 2000
rect 4098 1944 4660 1996
rect 4100 1930 4660 1944
rect 4740 1930 4750 2000
rect -1860 -1260 -1360 -1020
rect 2950 -1730 3140 -1660
rect 3130 -1780 3140 -1730
rect 3320 -1780 3330 -1660
rect 3140 -1810 3330 -1780
rect 3200 -2350 4620 -2270
rect -1390 -4120 -1380 -4020
rect -1270 -4120 -1260 -4020
rect 4180 -5090 4190 -5080
rect 4090 -5190 4190 -5090
rect 4180 -5200 4190 -5190
rect 4290 -5200 4300 -5080
rect 2840 -8140 2850 -7990
rect 3020 -8140 3030 -7990
rect 4470 -8030 4620 -2350
rect 3600 -8100 3650 -8030
rect 3790 -8100 3840 -8030
rect 3980 -8100 4030 -8030
rect 4170 -8100 4220 -8030
rect 4370 -8110 4420 -8040
rect 4560 -8110 4610 -8040
rect -1390 -8850 -1380 -8760
rect -1270 -8850 -1260 -8760
rect 3160 -8880 3570 -8800
rect 5060 -8880 5480 -8800
rect 5590 -8880 6130 -8810
rect 5390 -8910 5480 -8880
rect 5390 -9090 5440 -8910
rect 5500 -9090 5510 -8910
rect 5630 -9090 5640 -8910
rect 5700 -9090 5710 -8910
rect 5820 -9090 5830 -8910
rect 5890 -9090 5900 -8910
rect 5530 -9310 5540 -9150
rect 5600 -9310 5610 -9150
rect 5730 -9310 5740 -9150
rect 5800 -9310 5810 -9150
rect 5920 -9310 5930 -9150
rect 5990 -9310 6000 -9150
rect 6030 -9300 6130 -8880
rect 6030 -9340 6060 -9300
rect 3210 -9420 3500 -9340
rect 5480 -9410 6060 -9340
rect 6130 -9410 6140 -9300
rect 1330 -9890 6340 -9850
rect 1330 -9910 1380 -9890
rect 1210 -10040 1380 -9910
rect 1130 -10060 1380 -10040
rect 1330 -10960 1380 -10060
rect 6300 -10960 6340 -9890
rect 6380 -10070 6390 -9960
rect 6460 -10070 6470 -9960
rect 6390 -10130 6450 -10070
rect 6420 -10920 6480 -10140
rect 6664 -10200 6766 -10188
rect 6610 -10320 6620 -10200
rect 6760 -10320 6770 -10200
rect 6664 -10332 6766 -10320
rect 1330 -11010 6340 -10960
<< via1 >>
rect 4660 1930 4740 2000
rect 3140 -1780 3320 -1660
rect -1380 -4120 -1270 -4020
rect 4190 -5200 4290 -5080
rect 2850 -8140 3020 -7990
rect -1380 -8850 -1270 -8760
rect 5440 -9090 5500 -8910
rect 5640 -9090 5700 -8910
rect 5830 -9090 5890 -8910
rect 5540 -9310 5600 -9150
rect 5740 -9310 5800 -9150
rect 5930 -9310 5990 -9150
rect 6060 -9410 6130 -9300
rect 6390 -10070 6460 -9960
rect 6620 -10320 6670 -10200
rect 6670 -10320 6760 -10200
<< metal2 >>
rect 4660 2000 4740 2010
rect 4660 1920 4740 1930
rect 830 1750 1040 1890
rect 1800 670 1910 840
rect 1770 160 1890 320
rect 2720 -1460 2890 -1320
rect 3140 -1660 3320 -1650
rect 3140 -1790 3320 -1780
rect 1260 -2150 1530 -2140
rect 1260 -2430 1530 -2420
rect -1380 -4020 -1270 -4010
rect -1380 -8760 -1270 -4120
rect -1020 -4690 -910 -4530
rect 4190 -5080 4290 -5070
rect 5080 -5080 5170 -5070
rect 4290 -5200 5080 -5080
rect 4190 -5210 4290 -5200
rect 5080 -5210 5170 -5200
rect 3880 -5340 4500 -5260
rect 1700 -6390 1900 -6240
rect 1740 -6900 1920 -6760
rect 4320 -7540 4500 -5340
rect 4320 -7710 5050 -7540
rect 2850 -7990 3020 -7980
rect 2850 -8150 3020 -8140
rect 4550 -8090 4620 -8080
rect 4550 -8260 4620 -8250
rect 4930 -8540 5050 -7710
rect 2670 -8790 2920 -8600
rect 4930 -8650 6350 -8540
rect 4600 -8760 4720 -8660
rect -1380 -8860 -1270 -8850
rect 5440 -8910 5500 -8900
rect 5640 -8910 5700 -8900
rect 5830 -8910 5890 -8900
rect 5500 -9090 5640 -8910
rect 5700 -9090 5830 -8910
rect 5440 -9100 5500 -9090
rect 5640 -9100 5700 -9090
rect 5830 -9100 5890 -9090
rect 1250 -9210 1480 -9200
rect 3170 -9310 3550 -9140
rect 5540 -9150 5600 -9140
rect 5740 -9150 5800 -9140
rect 5930 -9150 5990 -9140
rect 5080 -9310 5540 -9150
rect 5600 -9310 5740 -9150
rect 5800 -9310 5930 -9150
rect 5540 -9320 5600 -9310
rect 5740 -9320 5800 -9310
rect 5930 -9320 5990 -9310
rect 6060 -9300 6130 -9290
rect 6060 -9420 6130 -9410
rect 1250 -9660 1480 -9650
rect 6230 -9700 6350 -8650
rect 6230 -9810 6760 -9700
rect 6390 -9960 6460 -9950
rect 6390 -10080 6460 -10070
rect 6620 -10200 6760 -9810
rect 6620 -10330 6760 -10320
<< via2 >>
rect 4660 1930 4740 2000
rect 3140 -1780 3320 -1660
rect 1260 -2420 1530 -2150
rect 5080 -5200 5170 -5080
rect 2850 -8140 3020 -7990
rect 4550 -8250 4620 -8090
rect 1250 -9650 1480 -9210
rect 6060 -9410 6130 -9300
rect 6390 -10070 6460 -9960
<< metal3 >>
rect 1040 1990 1140 2120
rect 4630 1910 4640 2020
rect 4760 1910 4770 2020
rect 2900 1040 3170 1170
rect 3130 -1660 3330 -1650
rect 3130 -1780 3140 -1660
rect 3320 -1780 3330 -1660
rect 3130 -2020 3330 -1780
rect 3140 -2140 3320 -2020
rect 1250 -2150 1540 -2145
rect 1250 -2420 1260 -2150
rect 1530 -2420 1540 -2150
rect 1250 -2425 1540 -2420
rect 630 -2970 700 -2870
rect 5070 -5080 5180 -5075
rect 5070 -5200 5080 -5080
rect 5170 -5200 5180 -5080
rect 5070 -5205 5180 -5200
rect 2920 -6050 3180 -5930
rect 2840 -7990 3030 -7985
rect 2840 -8140 2850 -7990
rect 3020 -8140 3030 -7990
rect 2840 -8145 3030 -8140
rect 4540 -8090 4630 -8085
rect 1240 -9210 1490 -9205
rect 2850 -9210 3020 -8145
rect 4540 -8250 4550 -8090
rect 4620 -8250 5190 -8090
rect 4540 -8255 4630 -8250
rect 1240 -9650 1250 -9210
rect 1480 -9650 1490 -9210
rect 6050 -9300 6140 -9295
rect 6050 -9410 6060 -9300
rect 6130 -9410 6460 -9300
rect 6050 -9415 6140 -9410
rect 1240 -9655 1490 -9650
rect 630 -10020 700 -9920
rect 6390 -9955 6460 -9410
rect 6380 -9960 6470 -9955
rect 6380 -10070 6390 -9960
rect 6460 -10070 6470 -9960
rect 6380 -10075 6470 -10070
<< via3 >>
rect 4640 2000 4760 2020
rect 4640 1930 4660 2000
rect 4660 1930 4740 2000
rect 4740 1930 4760 2000
rect 4640 1910 4760 1930
rect 1260 -2420 1530 -2150
rect 5080 -5200 5170 -5080
rect 1250 -9650 1480 -9210
<< metal4 >>
rect 4639 2020 4761 2021
rect 4639 1910 4640 2020
rect 4760 1960 4761 2020
rect 4760 1910 5080 1960
rect 4639 1909 5080 1910
rect 4640 1850 5080 1909
rect 1259 -2150 1531 -2149
rect 1259 -2260 1260 -2150
rect 1530 -2260 1531 -2150
rect 1530 -2420 2200 -2260
rect 1370 -2560 2200 -2420
rect 5060 -5080 5760 -4030
rect 5060 -5200 5080 -5080
rect 5170 -5200 5760 -5080
rect 5060 -5360 5760 -5200
rect 11390 -5310 11730 -4190
rect 1249 -9210 1481 -9209
rect 1249 -9380 1250 -9210
rect 1480 -9380 1481 -9210
rect 1480 -9650 1820 -9380
rect 1360 -9800 1820 -9650
<< via4 >>
rect 1090 -2420 1260 -2260
rect 1260 -2420 1370 -2260
rect 1090 -2560 1370 -2420
rect 1060 -9650 1250 -9380
rect 1250 -9650 1360 -9380
rect 1060 -9800 1360 -9650
<< metal5 >>
rect 3230 2360 5960 2680
rect 3230 1630 3590 2360
rect 5640 1880 5960 2360
rect 1066 -2260 1394 -2236
rect 1066 -2560 1090 -2260
rect 1370 -2560 1394 -2260
rect 1066 -2584 1394 -2560
rect 4360 -2680 5080 -2360
rect 5750 -4590 6070 -3980
rect 3300 -4970 6070 -4590
rect 3300 -5460 3680 -4970
rect 4680 -4980 6070 -4970
rect 5750 -5430 6070 -4980
rect 11110 -5520 11470 -3990
rect 1036 -9380 1384 -9356
rect 1036 -9800 1060 -9380
rect 1360 -9800 1384 -9380
rect 4300 -9750 5060 -9430
rect 1036 -9824 1384 -9800
use sky130_fd_pr__cap_mim_m3_1_J5CT7Z  sky130_fd_pr__cap_mim_m3_1_J5CT7Z_0
timestamp 1647254192
transform 1 0 3290 0 1 -10380
box -1650 -1300 1649 1300
use sky130_fd_pr__cap_mim_m3_1_J5CT7Z  sky130_fd_pr__cap_mim_m3_1_J5CT7Z_1
timestamp 1647254192
transform 1 0 3280 0 1 -3290
box -1650 -1300 1649 1300
use sky130_fd_pr__cap_mim_m3_2_LJ5JLG#0  sky130_fd_pr__cap_mim_m3_2_LJ5JLG_0
timestamp 1647254192
transform -1 0 8373 0 -1 -8409
box -3351 -3101 3373 3101
use sky130_fd_pr__cap_mim_m3_2_LJ5JLG#0  sky130_fd_pr__cap_mim_m3_2_LJ5JLG_1
timestamp 1647254192
transform -1 0 8373 0 -1 -1099
box -3351 -3101 3373 3101
use sky130_fd_pr__cap_var_lvt_MZUN4J  sky130_fd_pr__cap_var_lvt_MZUN4J_0
timestamp 1647254192
transform 1 0 3733 0 1 -10422
box -2283 -728 2283 728
use sky130_fd_pr__nfet_01v8_CDW43Z  sky130_fd_pr__nfet_01v8_CDW43Z_0
timestamp 1647254192
transform 1 0 6476 0 1 -10820
box -296 -260 296 260
use sky130_fd_pr__nfet_01v8_SC2JGL  sky130_fd_pr__nfet_01v8_SC2JGL_0
timestamp 1647254192
transform 1 0 5717 0 1 -9110
box -407 -410 407 410
use sky130_fd_pr__pfet_01v8_GCYTE7  sky130_fd_pr__pfet_01v8_GCYTE7_0
timestamp 1647254192
transform 1 0 6476 0 1 -10261
box -296 -269 296 269
use tia_cur_mirror  tia_cur_mirror_0
timestamp 1647254192
transform 1 0 3420 0 1 -8620
box -60 -900 1822 740
use tia_one_tia  tia_one_tia_0
timestamp 1647269090
transform 1 0 614 0 1 -890
box -2010 -3360 3840 3680
use tia_one_tia  tia_one_tia_1
timestamp 1647269090
transform 1 0 614 0 1 -7960
box -2010 -3360 3840 3680
<< labels >>
rlabel metal1 -1840 -1240 -1560 -1040 1 Input
port 6 n
rlabel metal4 11480 -4560 11690 -4360 1 VN
port 8 n
rlabel metal2 2720 -1460 2890 -1320 3 VM5D
rlabel metal3 1040 1990 1140 2120 1 Out_1
port 4 n
rlabel metal2 4600 -8760 4720 -8660 1 VM6D
rlabel metal3 6390 -9510 6450 -9410 1 Disable_TIA
port 5 n
rlabel metal1 6090 -9890 6150 -9850 1 Disable_TIA_B
rlabel metal3 630 -10020 700 -9920 1 VM40D
rlabel metal3 630 -2970 700 -2870 1 VM28D
rlabel metal3 5080 -8250 5190 -8090 1 I_Bias1
port 7 n
rlabel metal2 1800 670 1910 840 1 Out_1
rlabel metal3 2900 1040 3170 1170 1 Out_2
port 2 n
rlabel metal5 11130 -5060 11230 -4890 1 VPP
port 1 n
rlabel metal3 2920 -6050 3180 -5930 1 VM31D
rlabel metal2 1700 -6390 1900 -6240 1 Out_ref
rlabel metal2 1740 -6900 1920 -6760 1 VM39D
rlabel metal2 2670 -8790 2920 -8600 1 VM36D
<< end >>
