magic
tech sky130A
magscale 1 2
timestamp 1647254192
<< pwell >>
rect -1367 -1598 1367 1598
<< psubdiff >>
rect -1331 1528 -1235 1562
rect 1235 1528 1331 1562
rect -1331 1466 -1297 1528
rect 1297 1466 1331 1528
rect -1331 -1528 -1297 -1466
rect 1297 -1528 1331 -1466
rect -1331 -1562 -1235 -1528
rect 1235 -1562 1331 -1528
<< psubdiffcont >>
rect -1235 1528 1235 1562
rect -1331 -1466 -1297 1466
rect 1297 -1466 1331 1466
rect -1235 -1562 1235 -1528
<< xpolycontact >>
rect -1201 1000 -919 1432
rect -1201 -1432 -919 -1000
rect -671 1000 -389 1432
rect -671 -1432 -389 -1000
rect -141 1000 141 1432
rect -141 -1432 141 -1000
rect 389 1000 671 1432
rect 389 -1432 671 -1000
rect 919 1000 1201 1432
rect 919 -1432 1201 -1000
<< xpolyres >>
rect -1201 -1000 -919 1000
rect -671 -1000 -389 1000
rect -141 -1000 141 1000
rect 389 -1000 671 1000
rect 919 -1000 1201 1000
<< locali >>
rect -1331 1528 -1235 1562
rect 1235 1528 1331 1562
rect -1331 1466 -1297 1528
rect 1297 1466 1331 1528
rect -1331 -1528 -1297 -1466
rect 1297 -1528 1331 -1466
rect -1331 -1562 -1235 -1528
rect 1235 -1562 1331 -1528
<< viali >>
rect -1185 1017 -935 1414
rect -655 1017 -405 1414
rect -125 1017 125 1414
rect 405 1017 655 1414
rect 935 1017 1185 1414
rect -1185 -1414 -935 -1017
rect -655 -1414 -405 -1017
rect -125 -1414 125 -1017
rect 405 -1414 655 -1017
rect 935 -1414 1185 -1017
<< metal1 >>
rect -1191 1414 -929 1426
rect -1191 1017 -1185 1414
rect -935 1017 -929 1414
rect -1191 1005 -929 1017
rect -661 1414 -399 1426
rect -661 1017 -655 1414
rect -405 1017 -399 1414
rect -661 1005 -399 1017
rect -131 1414 131 1426
rect -131 1017 -125 1414
rect 125 1017 131 1414
rect -131 1005 131 1017
rect 399 1414 661 1426
rect 399 1017 405 1414
rect 655 1017 661 1414
rect 399 1005 661 1017
rect 929 1414 1191 1426
rect 929 1017 935 1414
rect 1185 1017 1191 1414
rect 929 1005 1191 1017
rect -1191 -1017 -929 -1005
rect -1191 -1414 -1185 -1017
rect -935 -1414 -929 -1017
rect -1191 -1426 -929 -1414
rect -661 -1017 -399 -1005
rect -661 -1414 -655 -1017
rect -405 -1414 -399 -1017
rect -661 -1426 -399 -1414
rect -131 -1017 131 -1005
rect -131 -1414 -125 -1017
rect 125 -1414 131 -1017
rect -131 -1426 131 -1414
rect 399 -1017 661 -1005
rect 399 -1414 405 -1017
rect 655 -1414 661 -1017
rect 399 -1426 661 -1414
rect 929 -1017 1191 -1005
rect 929 -1414 935 -1017
rect 1185 -1414 1191 -1017
rect 929 -1426 1191 -1414
<< res1p41 >>
rect -1203 -1002 -917 1002
rect -673 -1002 -387 1002
rect -143 -1002 143 1002
rect 387 -1002 673 1002
rect 917 -1002 1203 1002
<< properties >>
string FIXED_BBOX -1314 -1545 1314 1545
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 10 m 1 nx 5 wmin 1.410 lmin 0.50 rho 2000 val 14.451k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
