magic
tech sky130A
magscale 1 2
timestamp 1646921651
<< error_p >>
rect -125 272 -67 278
rect 67 272 125 278
rect -125 238 -113 272
rect 67 238 79 272
rect -125 232 -67 238
rect 67 232 125 238
rect -221 -238 -163 -232
rect -29 -238 29 -232
rect 163 -238 221 -232
rect -221 -272 -209 -238
rect -29 -272 -17 -238
rect 163 -272 175 -238
rect -221 -278 -163 -272
rect -29 -278 29 -272
rect 163 -278 221 -272
<< pwell >>
rect -407 -410 407 410
<< nmos >>
rect -207 -200 -177 200
rect -111 -200 -81 200
rect -15 -200 15 200
rect 81 -200 111 200
rect 177 -200 207 200
<< ndiff >>
rect -269 188 -207 200
rect -269 -188 -257 188
rect -223 -188 -207 188
rect -269 -200 -207 -188
rect -177 188 -111 200
rect -177 -188 -161 188
rect -127 -188 -111 188
rect -177 -200 -111 -188
rect -81 188 -15 200
rect -81 -188 -65 188
rect -31 -188 -15 188
rect -81 -200 -15 -188
rect 15 188 81 200
rect 15 -188 31 188
rect 65 -188 81 188
rect 15 -200 81 -188
rect 111 188 177 200
rect 111 -188 127 188
rect 161 -188 177 188
rect 111 -200 177 -188
rect 207 188 269 200
rect 207 -188 223 188
rect 257 -188 269 188
rect 207 -200 269 -188
<< ndiffc >>
rect -257 -188 -223 188
rect -161 -188 -127 188
rect -65 -188 -31 188
rect 31 -188 65 188
rect 127 -188 161 188
rect 223 -188 257 188
<< psubdiff >>
rect -371 340 -275 374
rect 275 340 371 374
rect -371 278 -337 340
rect 337 278 371 340
rect -371 -340 -337 -278
rect 337 -340 371 -278
rect -371 -374 -275 -340
rect 275 -374 371 -340
<< psubdiffcont >>
rect -275 340 275 374
rect -371 -278 -337 278
rect 337 -278 371 278
rect -275 -374 275 -340
<< poly >>
rect -129 272 -63 288
rect -129 238 -113 272
rect -79 238 -63 272
rect -207 200 -177 226
rect -129 222 -63 238
rect 63 272 129 288
rect 63 238 79 272
rect 113 238 129 272
rect -111 200 -81 222
rect -15 200 15 226
rect 63 222 129 238
rect 81 200 111 222
rect 177 200 207 226
rect -207 -222 -177 -200
rect -225 -238 -159 -222
rect -111 -226 -81 -200
rect -15 -222 15 -200
rect -225 -272 -209 -238
rect -175 -272 -159 -238
rect -225 -288 -159 -272
rect -33 -238 33 -222
rect 81 -226 111 -200
rect 177 -222 207 -200
rect -33 -272 -17 -238
rect 17 -272 33 -238
rect -33 -288 33 -272
rect 159 -238 225 -222
rect 159 -272 175 -238
rect 209 -272 225 -238
rect 159 -288 225 -272
<< polycont >>
rect -113 238 -79 272
rect 79 238 113 272
rect -209 -272 -175 -238
rect -17 -272 17 -238
rect 175 -272 209 -238
<< locali >>
rect -371 340 -275 374
rect 275 340 371 374
rect -371 278 -337 340
rect 337 278 371 340
rect -129 238 -113 272
rect -79 238 -63 272
rect 63 238 79 272
rect 113 238 129 272
rect -257 188 -223 204
rect -257 -204 -223 -188
rect -161 188 -127 204
rect -161 -204 -127 -188
rect -65 188 -31 204
rect -65 -204 -31 -188
rect 31 188 65 204
rect 31 -204 65 -188
rect 127 188 161 204
rect 127 -204 161 -188
rect 223 188 257 204
rect 223 -204 257 -188
rect -225 -272 -209 -238
rect -175 -272 -159 -238
rect -33 -272 -17 -238
rect 17 -272 33 -238
rect 159 -272 175 -238
rect 209 -272 225 -238
rect -371 -340 -337 -278
rect 337 -340 371 -278
rect -371 -374 -275 -340
rect 275 -374 371 -340
<< viali >>
rect -113 238 -79 272
rect 79 238 113 272
rect -257 -188 -223 188
rect -161 -188 -127 188
rect -65 -188 -31 188
rect 31 -188 65 188
rect 127 -188 161 188
rect 223 -188 257 188
rect -209 -272 -175 -238
rect -17 -272 17 -238
rect 175 -272 209 -238
<< metal1 >>
rect -125 272 -67 278
rect -125 238 -113 272
rect -79 238 -67 272
rect -125 232 -67 238
rect 67 272 125 278
rect 67 238 79 272
rect 113 238 125 272
rect 67 232 125 238
rect -263 188 -217 200
rect -263 -188 -257 188
rect -223 -188 -217 188
rect -263 -200 -217 -188
rect -167 188 -121 200
rect -167 -188 -161 188
rect -127 -188 -121 188
rect -167 -200 -121 -188
rect -71 188 -25 200
rect -71 -188 -65 188
rect -31 -188 -25 188
rect -71 -200 -25 -188
rect 25 188 71 200
rect 25 -188 31 188
rect 65 -188 71 188
rect 25 -200 71 -188
rect 121 188 167 200
rect 121 -188 127 188
rect 161 -188 167 188
rect 121 -200 167 -188
rect 217 188 263 200
rect 217 -188 223 188
rect 257 -188 263 188
rect 217 -200 263 -188
rect -221 -238 -163 -232
rect -221 -272 -209 -238
rect -175 -272 -163 -238
rect -221 -278 -163 -272
rect -29 -238 29 -232
rect -29 -272 -17 -238
rect 17 -272 29 -238
rect -29 -278 29 -272
rect 163 -238 221 -232
rect 163 -272 175 -238
rect 209 -272 221 -238
rect 163 -278 221 -272
<< properties >>
string FIXED_BBOX -354 -357 354 357
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.150 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
