* NGSPICE file created from tia_core_flat.ext - technology: sky130A

.subckt tia_core_flat Out_2 Out_1 Disable_TIA I_Bias1 Input VN VPP
X0 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=6.432e+13p pd=4.8032e+08u as=3.412e+13p ps=2.6612e+08u w=2e+06u l=200000u
X1 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=6.432e+13p pd=4.8032e+08u as=3.412e+13p ps=2.6612e+08u w=2e+06u l=200000u
X2 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X3 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X4 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X5 Out_2 Out_1 Input Input sky130_fd_pr__nfet_01v8_lvt ad=9.28e+12p pd=7.328e+07u as=9.28e+12p ps=7.328e+07u w=2e+06u l=200000u
X6 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=1.01615e+14p pd=6.645e+08u as=0p ps=0u w=2e+06u l=150000u
X7 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8 w_2300_n7574# a_n1188_n8454# a_2412_n5577# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=9.28e+12p pd=7.328e+07u as=9.28e+12p ps=7.328e+07u w=2e+06u l=200000u
X9 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=4.3065e+13p pd=3.405e+08u as=1.856e+13p ps=1.4656e+08u w=2e+06u l=200000u
X10 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X11 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X14 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X16 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X17 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X18 w_2300_n7574# a_n1188_n8454# a_2412_n5577# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X19 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X20 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X21 a_2412_n5577# a_n1188_n8454# w_2300_n7574# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X22 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X23 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X24 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=1.856e+13p pd=1.4656e+08u as=0p ps=0u w=2e+06u l=200000u
X25 VM5D I_Bias1 Out_1 VN sky130_fd_pr__nfet_01v8 ad=6.28e+12p pd=4.628e+07u as=0p ps=0u w=2e+06u l=150000u
X26 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X27 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X28 VPP VN Out_2 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+12p ps=2.748e+07u w=2e+06u l=500000u
X29 Out_2 Out_1 Input Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X30 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X31 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X32 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X33 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X34 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X35 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X36 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X37 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X38 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X39 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X40 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X41 a_n1188_n8454# I_Bias1 a_1602_n8490# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.28e+12p ps=4.628e+07u w=2e+06u l=150000u
X42 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X43 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X44 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X45 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X46 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X47 w_2300_n7574# a_n1188_n8454# a_2412_n5577# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X48 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X49 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X50 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X51 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X52 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X53 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X54 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X55 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X56 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X57 VPP VN sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X58 w_2300_n7574# a_n1188_n8454# a_2412_n5577# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X59 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X60 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X61 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X62 a_1602_n8490# I_Bias1 a_n1188_n8454# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X63 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X64 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X65 a_2412_n5577# a_n1188_n8454# w_2300_n7574# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X66 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X67 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X68 VN I_Bias1 VM6D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.28e+12p ps=4.628e+07u w=2e+06u l=1e+06u
X69 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X70 Out_1 I_Bias1 VM5D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X71 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X72 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X73 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X74 a_2412_n5577# a_n1188_n8454# w_2300_n7574# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X75 VN I_Bias1 a_1602_n8490# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X76 a_n1188_n8454# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X77 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X78 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X79 a_n1188_n8454# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X80 Out_1 I_Bias1 VM5D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X81 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X82 a_n1188_n8454# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X83 Out_2 Out_1 Input Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X84 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X85 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X86 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X87 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X88 VPP Disable_TIA Disable_TIA_B VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.45e+11p ps=1.58e+06u w=500000u l=1e+06u
X89 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X90 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X91 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X92 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X93 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X94 Out_2 Out_1 Input Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X95 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X96 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X97 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X98 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X99 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X100 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X101 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X102 VPP VN Out_2 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X103 a_1602_n8490# I_Bias1 a_n1188_n8454# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X104 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X105 w_2300_n7574# a_n1188_n8454# a_2412_n5577# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X106 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X107 a_1602_n8490# I_Bias1 VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X108 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X109 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X110 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X111 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X112 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X113 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X114 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X115 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X116 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X117 w_2300_n7574# a_n1188_n8454# a_2412_n5577# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X118 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X119 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X120 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X121 a_n1188_n8454# I_Bias1 a_1602_n8490# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X122 w_2300_n7574# a_n1188_n8454# a_2412_n5577# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X123 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X124 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X125 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X126 VM5D I_Bias1 VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X127 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X128 a_n1188_n8454# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X129 a_n1188_n8454# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X130 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X131 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X132 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X133 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X134 VM5D I_Bias1 Out_1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X135 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X136 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X137 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X138 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X139 a_n1188_n8454# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X140 a_n1188_n8454# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X141 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X142 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X143 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X144 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X145 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X146 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X147 I_Bias1 I_Bias1 VM6D VN sky130_fd_pr__nfet_01v8 ad=5.9e+12p pd=4.19e+07u as=0p ps=0u w=2e+06u l=150000u
X148 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X149 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X150 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X151 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X152 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X153 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X154 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X155 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X156 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X157 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X158 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X159 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X160 VPP VN Out_2 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X161 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X162 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X163 a_n1188_n8454# I_Bias1 a_1602_n8490# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X164 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X165 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X166 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X167 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X168 VPP VN a_2412_n5577# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+12p ps=2.748e+07u w=2e+06u l=500000u
X169 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X170 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X171 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X172 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X173 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X174 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X175 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X176 a_n1188_n8454# I_Bias1 a_1602_n8490# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X177 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X178 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X179 VN I_Bias1 sky130_fd_pr__cap_mim_m3_1 l=1.2e+07u w=1.5e+07u
X180 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X181 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X182 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X183 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X184 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X185 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X186 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X187 a_2412_n5577# a_n1188_n8454# w_2300_n7574# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X188 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X189 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X190 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X191 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X192 VPP VN a_2412_n5577# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X193 a_n1188_n8454# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X194 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X195 Out_2 Out_1 Input Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X196 a_2412_n5577# a_n1188_n8454# w_2300_n7574# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X197 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X198 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X199 a_1602_n8490# I_Bias1 a_n1188_n8454# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X200 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X201 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X202 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X203 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X204 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X205 VM6D I_Bias1 I_Bias1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X206 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X207 a_n1188_n8454# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X208 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X209 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X210 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X211 VM6D I_Bias1 VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X212 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X213 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X214 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X215 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X216 Out_2 Out_1 Input Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X217 VN Disable_TIA Disable_TIA_B VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.45e+11p ps=1.58e+06u w=500000u l=1e+06u
X218 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X219 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X220 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X221 a_n1188_n8454# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X222 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X223 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X224 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X225 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X226 a_2412_n5577# VN VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X227 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X228 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X229 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X230 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X231 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X232 VM6D I_Bias1 I_Bias1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X233 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X234 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X235 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X236 w_2300_n7574# a_n1188_n8454# a_2412_n5577# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X237 a_2412_n5577# VN VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X238 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X239 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X240 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X241 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X242 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X243 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X244 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X245 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X246 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X247 a_1602_n8490# I_Bias1 a_n1188_n8454# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X248 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X249 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X250 VN I_Bias1 VM5D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X251 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X252 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X253 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X254 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X255 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X256 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X257 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X258 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X259 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X260 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X261 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X262 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X263 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X264 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X265 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X266 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X267 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X268 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X269 VN Disable_TIA I_Bias1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X270 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X271 VN I_Bias1 sky130_fd_pr__cap_mim_m3_1 l=1.2e+07u w=1.5e+07u
X272 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X273 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X274 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X275 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X276 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X277 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X278 VM6D I_Bias1 I_Bias1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X279 a_2412_n5577# a_n1188_n8454# w_2300_n7574# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X280 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X281 Out_2 Out_1 Input Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X282 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X283 I_Bias1 I_Bias1 VM6D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X284 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X285 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X286 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X287 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X288 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X289 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X290 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X291 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X292 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X293 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X294 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X295 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X296 I_Bias1 I_Bias1 VM6D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X297 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X298 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X299 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X300 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X301 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X302 Out_2 Out_1 Input Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X303 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X304 a_n1188_n8454# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X305 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X306 a_n1188_n8454# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X307 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X308 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X309 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X310 Out_1 I_Bias1 VM5D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X311 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X312 VM5D I_Bias1 VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X313 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X314 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X315 w_2300_n7574# a_n1188_n8454# a_2412_n5577# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X316 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X317 VPP VN Out_2 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X318 a_n1188_n8454# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X319 a_n1188_n8454# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X320 Out_2 VN VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X321 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X322 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X323 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X324 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X325 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X326 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X327 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X328 w_2300_n7574# a_n1188_n8454# a_2412_n5577# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X329 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X330 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X331 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X332 VM5D I_Bias1 Out_1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X333 I_Bias1 I_Bias1 VM6D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X334 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X335 a_2412_n5577# a_n1188_n8454# w_2300_n7574# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X336 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X337 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X338 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X339 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X340 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X341 VN I_Bias1 VM5D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X342 Out_2 VN VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X343 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X344 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X345 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X346 a_2412_n5577# a_n1188_n8454# w_2300_n7574# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X347 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X348 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X349 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X350 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X351 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X352 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X353 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X354 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X355 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X356 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X357 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X358 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X359 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X360 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X361 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X362 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X363 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X364 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X365 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X366 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X367 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X368 VM5D I_Bias1 Out_1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X369 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X370 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X371 a_1602_n8490# I_Bias1 VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X372 a_2412_n5577# a_n1188_n8454# w_2300_n7574# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X373 VPP VN sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X374 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X375 Out_2 Out_1 Input Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X376 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X377 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X378 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X379 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X380 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X381 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X382 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X383 a_2412_n5577# a_n1188_n8454# w_2300_n7574# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X384 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X385 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X386 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X387 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X388 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X389 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X390 Out_1 I_Bias1 VM5D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X391 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X392 a_n1188_n8454# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X393 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X394 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X395 Out_2 Out_1 Input Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X396 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X397 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X398 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X399 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X400 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X401 VPP VN a_2412_n5577# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X402 a_n1188_n8454# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X403 w_2300_n7574# a_n1188_n8454# a_2412_n5577# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X404 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X405 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X406 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X407 VN I_Bias1 VM6D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X408 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X409 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X410 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X411 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X412 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X413 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X414 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X415 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X416 w_2300_n7574# a_n1188_n8454# a_2412_n5577# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X417 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X418 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X419 a_1602_n8490# I_Bias1 a_n1188_n8454# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X420 Out_2 VN VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X421 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X422 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X423 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X424 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X425 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X426 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X427 Out_1 I_Bias1 VM5D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X428 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X429 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X430 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X431 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X432 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X433 a_2412_n5577# VN VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X434 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X435 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X436 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X437 VM6D I_Bias1 VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X438 Out_1 I_Bias1 VM5D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X439 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X440 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X441 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X442 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X443 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X444 a_2412_n5577# a_n1188_n8454# w_2300_n7574# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X445 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X446 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X447 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X448 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X449 a_2412_n5577# a_n1188_n8454# w_2300_n7574# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X450 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X451 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X452 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X453 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X454 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X455 Disable_TIA_B VN VN sky130_fd_pr__cap_var_lvt pd=0u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X456 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X457 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X458 VM5D I_Bias1 Out_1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X459 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X460 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X461 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X462 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X463 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X464 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X465 a_n1188_n8454# I_Bias1 a_1602_n8490# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X466 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X467 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X468 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X469 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X470 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X471 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X472 Out_2 Out_1 Input Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X473 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X474 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X475 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X476 VN I_Bias1 a_1602_n8490# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X477 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X478 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X479 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X480 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X481 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X482 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X483 VPP VN a_2412_n5577# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X484 a_n1188_n8454# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X485 a_n1188_n8454# I_Bias1 a_1602_n8490# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X486 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X487 w_2300_n7574# a_n1188_n8454# a_2412_n5577# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X488 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X489 Disable_TIA_B VN VN sky130_fd_pr__cap_var_lvt pd=0u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X490 a_n1188_n8454# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X491 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X492 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X493 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X494 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X495 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X496 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X497 I_Bias1 Disable_TIA VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X498 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X499 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X500 a_n1188_n8454# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X501 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X502 VM5D I_Bias1 Out_1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X503 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X504 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X505 VN I_Bias1 VM5D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X506 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X507 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X508 Disable_TIA_B VN VN sky130_fd_pr__cap_var_lvt pd=0u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X509 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X510 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X511 I_Bias1 I_Bias1 VM6D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X512 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X513 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X514 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X515 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X516 Out_2 VN VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X517 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X518 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X519 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X520 w_2300_n7574# a_n1188_n8454# a_2412_n5577# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X521 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X522 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X523 Disable_TIA_B VN VN sky130_fd_pr__cap_var_lvt pd=0u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X524 a_2412_n5577# VN VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X525 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X526 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X527 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X528 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X529 VPP m4_n1346_n2030# sky130_fd_pr__cap_mim_m3_2 l=1.8e+07u w=2.5e+07u
X530 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X531 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X532 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X533 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X534 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X535 w_2300_n7574# a_n1188_n8454# a_2412_n5577# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X536 VM6D I_Bias1 I_Bias1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X537 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X538 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X539 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X540 w_2300_n7574# a_n1188_n8454# a_2412_n5577# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X541 VM6D I_Bias1 VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X542 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X543 VM5D I_Bias1 VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X544 VPP VN Out_2 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X545 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X546 a_1602_n8490# I_Bias1 a_n1188_n8454# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X547 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X548 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X549 a_n1188_n8454# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X550 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X551 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X552 a_1602_n8490# I_Bias1 VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X553 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X554 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X555 Disable_TIA_B VN VN sky130_fd_pr__cap_var_lvt pd=0u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X556 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X557 a_n1188_n8454# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X558 a_n1188_n8454# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X559 a_n1188_n8454# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X560 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X561 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X562 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X563 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X564 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X565 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X566 VM6D I_Bias1 I_Bias1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X567 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X568 VN Disable_TIA I_Bias1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X569 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X570 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X571 a_n1188_n8454# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X572 a_n1188_n8454# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X573 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X574 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X575 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X576 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X577 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X578 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X579 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X580 VN I_Bias1 a_1602_n8490# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X581 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X582 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X583 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X584 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X585 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X586 I_Bias1 Disable_TIA VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X587 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X588 VM6D I_Bias1 I_Bias1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X589 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X590 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X591 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X592 VPP m4_n1346_n9100# sky130_fd_pr__cap_mim_m3_2 l=1.8e+07u w=2.5e+07u
X593 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X594 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X595 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X596 Out_2 Out_1 Input Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X597 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X598 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X599 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X600 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X601 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X602 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X603 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X604 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X605 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X606 a_2412_n5577# VN VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X607 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X608 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X609 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X610 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X611 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X612 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X613 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X614 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X615 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X616 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X617 Out_2 Out_1 Input Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X618 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X619 a_n1188_n8454# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X620 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X621 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X622 Input Out_1 Out_2 Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X623 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X624 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X625 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X626 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X627 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X628 a_n1188_n8454# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X629 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X630 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X631 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X632 VN Disable_TIA_B VM40D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X633 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X634 a_n1188_n8454# w_2300_n7574# VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X635 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X636 Out_2 VN VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X637 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X638 VPP VN a_2412_n5577# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X639 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X640 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X641 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X642 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X643 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X644 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X645 a_n1188_n8454# w_2300_n7574# VM40D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X646 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X647 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X648 Out_2 Out_1 Input Input sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X649 I_Bias1 I_Bias1 VM6D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X650 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X651 VN Disable_TIA_B VM28D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X652 a_2412_n5577# a_n1188_n8454# w_2300_n7574# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X653 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X654 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X655 Out_1 Input VPP VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X656 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X657 VN I_Bias1 VM6D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X658 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X659 VPP Input Out_1 VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X660 Out_1 Input VM28D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X661 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X662 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X663 VM28D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X664 a_2412_n5577# a_n1188_n8454# w_2300_n7574# w_2300_n7574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X665 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X666 VPP w_2300_n7574# a_n1188_n8454# VPP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X667 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X668 VN Disable_TIA I_Bias1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X669 VM28D Input Out_1 VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X670 VM40D w_2300_n7574# a_n1188_n8454# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X671 VM40D Disable_TIA_B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

