magic
tech sky130A
magscale 1 2
timestamp 1646921651
<< locali >>
rect -30 3380 500 3450
rect -30 2690 40 3380
rect 430 2690 500 3380
rect -30 2600 820 2690
rect -30 2580 40 2600
rect 460 2580 820 2600
rect -30 40 130 2580
rect 660 40 820 2580
rect -30 -30 820 40
<< metal1 >>
rect 250 3270 470 3340
rect 198 3080 208 3240
rect 262 3080 272 3240
rect 100 2840 110 3000
rect 164 2840 174 3000
rect 296 2840 306 3000
rect 360 2840 370 3000
rect 398 2810 470 3270
rect 140 2740 470 2810
rect 230 2520 300 2740
rect 150 2470 630 2520
rect 100 2034 110 2194
rect 164 2034 174 2194
rect 230 2000 300 2470
rect 358 2274 368 2434
rect 422 2274 432 2434
rect 616 2034 626 2194
rect 680 2034 690 2194
rect 150 1850 630 2000
rect 100 1416 110 1576
rect 164 1416 174 1576
rect 230 1380 300 1850
rect 358 1656 368 1816
rect 422 1656 432 1816
rect 616 1416 626 1576
rect 680 1416 690 1576
rect 150 1230 630 1380
rect 100 1038 110 1198
rect 164 1038 174 1198
rect 230 770 300 1230
rect 616 1038 626 1198
rect 680 1038 690 1198
rect 358 798 368 958
rect 422 798 432 958
rect 150 610 630 770
rect 100 180 110 340
rect 164 180 174 340
rect 230 150 300 610
rect 358 420 368 580
rect 422 420 432 580
rect 616 180 626 340
rect 680 180 690 340
rect 150 90 630 150
<< via1 >>
rect 208 3080 262 3240
rect 110 2840 164 3000
rect 306 2840 360 3000
rect 110 2034 164 2194
rect 368 2274 422 2434
rect 626 2034 680 2194
rect 110 1416 164 1576
rect 368 1656 422 1816
rect 626 1416 680 1576
rect 110 1038 164 1198
rect 626 1038 680 1198
rect 368 798 422 958
rect 110 180 164 340
rect 368 420 422 580
rect 626 180 680 340
<< metal2 >>
rect 208 3240 262 3250
rect 208 3070 262 3080
rect 110 3000 530 3010
rect 164 2840 306 3000
rect 360 2840 530 3000
rect 110 2830 530 2840
rect 270 2434 530 2830
rect 270 2274 368 2434
rect 422 2274 530 2434
rect 10 2194 200 2210
rect 10 2034 110 2194
rect 164 2034 200 2194
rect 10 1576 200 2034
rect 10 1416 110 1576
rect 164 1416 200 1576
rect 10 1198 200 1416
rect 10 1038 110 1198
rect 164 1038 200 1198
rect 10 340 200 1038
rect 270 1816 530 2274
rect 270 1656 368 1816
rect 422 1656 530 1816
rect 270 958 530 1656
rect 270 798 368 958
rect 422 798 530 958
rect 270 580 530 798
rect 270 420 368 580
rect 422 420 530 580
rect 270 410 530 420
rect 580 2194 770 2210
rect 580 2034 626 2194
rect 680 2034 770 2194
rect 580 1576 770 2034
rect 580 1416 626 1576
rect 680 1416 770 1576
rect 580 1198 770 1416
rect 580 1038 626 1198
rect 680 1038 770 1198
rect 580 340 770 1038
rect 10 180 110 340
rect 164 180 626 340
rect 680 180 770 340
rect 10 -30 770 180
use sky130_fd_pr__nfet_01v8_M8466X  sky130_fd_pr__nfet_01v8_M8466X_0
timestamp 1646921651
transform 1 0 395 0 1 1307
box -425 -1337 425 1337
use sky130_fd_pr__nfet_01v8_WS53KN  sky130_fd_pr__nfet_01v8_WS53KN_0
timestamp 1646921651
transform 1 0 235 0 1 3040
box -265 -410 265 410
<< end >>
