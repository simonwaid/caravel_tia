magic
tech sky130A
magscale 1 2
timestamp 1647254192
<< poly >>
rect 182 9230 1208 9246
rect 182 9196 294 9230
rect 328 9196 486 9230
rect 520 9196 678 9230
rect 712 9196 870 9230
rect 904 9196 1062 9230
rect 1096 9196 1208 9230
rect 182 9180 1208 9196
rect 1560 9230 2586 9246
rect 1560 9196 1672 9230
rect 1706 9196 1864 9230
rect 1898 9196 2056 9230
rect 2090 9196 2248 9230
rect 2282 9196 2440 9230
rect 2474 9196 2586 9230
rect 1560 9180 2586 9196
rect 182 8720 1208 8736
rect 182 8686 198 8720
rect 232 8686 390 8720
rect 424 8686 582 8720
rect 616 8686 774 8720
rect 808 8686 966 8720
rect 1000 8686 1158 8720
rect 1192 8686 1208 8720
rect 182 8670 1208 8686
rect 1560 8720 2586 8736
rect 1560 8686 1576 8720
rect 1610 8686 1768 8720
rect 1802 8686 1960 8720
rect 1994 8686 2152 8720
rect 2186 8686 2344 8720
rect 2378 8686 2536 8720
rect 2570 8686 2586 8720
rect 1560 8670 2586 8686
rect 182 8612 1208 8628
rect 182 8578 198 8612
rect 232 8578 390 8612
rect 424 8578 582 8612
rect 616 8578 774 8612
rect 808 8578 966 8612
rect 1000 8578 1158 8612
rect 1192 8578 1208 8612
rect 182 8562 1208 8578
rect 1560 8612 2586 8628
rect 1560 8578 1576 8612
rect 1610 8578 1768 8612
rect 1802 8578 1960 8612
rect 1994 8578 2152 8612
rect 2186 8578 2344 8612
rect 2378 8578 2536 8612
rect 2570 8578 2586 8612
rect 1560 8562 2586 8578
rect 182 8102 1208 8118
rect 182 8068 296 8102
rect 330 8068 486 8102
rect 520 8068 678 8102
rect 712 8068 870 8102
rect 904 8068 1062 8102
rect 1096 8068 1208 8102
rect 182 8052 1208 8068
rect 1560 8102 2586 8118
rect 1560 8068 1672 8102
rect 1706 8068 1864 8102
rect 1898 8068 2056 8102
rect 2090 8068 2248 8102
rect 2282 8068 2438 8102
rect 2472 8068 2586 8102
rect 1560 8052 2586 8068
<< polycont >>
rect 294 9196 328 9230
rect 486 9196 520 9230
rect 678 9196 712 9230
rect 870 9196 904 9230
rect 1062 9196 1096 9230
rect 1672 9196 1706 9230
rect 1864 9196 1898 9230
rect 2056 9196 2090 9230
rect 2248 9196 2282 9230
rect 2440 9196 2474 9230
rect 198 8686 232 8720
rect 390 8686 424 8720
rect 582 8686 616 8720
rect 774 8686 808 8720
rect 966 8686 1000 8720
rect 1158 8686 1192 8720
rect 1576 8686 1610 8720
rect 1768 8686 1802 8720
rect 1960 8686 1994 8720
rect 2152 8686 2186 8720
rect 2344 8686 2378 8720
rect 2536 8686 2570 8720
rect 198 8578 232 8612
rect 390 8578 424 8612
rect 582 8578 616 8612
rect 774 8578 808 8612
rect 966 8578 1000 8612
rect 1158 8578 1192 8612
rect 1576 8578 1610 8612
rect 1768 8578 1802 8612
rect 1960 8578 1994 8612
rect 2152 8578 2186 8612
rect 2344 8578 2378 8612
rect 2536 8578 2570 8612
rect 296 8068 330 8102
rect 486 8068 520 8102
rect 678 8068 712 8102
rect 870 8068 904 8102
rect 1062 8068 1096 8102
rect 1672 8068 1706 8102
rect 1864 8068 1898 8102
rect 2056 8068 2090 8102
rect 2248 8068 2282 8102
rect 2438 8068 2472 8102
<< locali >>
rect 182 9196 294 9230
rect 328 9196 486 9230
rect 520 9196 678 9230
rect 712 9196 870 9230
rect 904 9196 1062 9230
rect 1096 9196 1208 9230
rect 1560 9196 1672 9230
rect 1706 9196 1864 9230
rect 1898 9196 2056 9230
rect 2090 9196 2248 9230
rect 2282 9196 2440 9230
rect 2474 9196 2586 9230
rect 182 8686 198 8720
rect 232 8686 390 8720
rect 424 8686 582 8720
rect 616 8686 774 8720
rect 808 8686 966 8720
rect 1000 8686 1158 8720
rect 1192 8686 1208 8720
rect 1560 8686 1576 8720
rect 1610 8686 1768 8720
rect 1802 8686 1960 8720
rect 1994 8686 2152 8720
rect 2186 8686 2344 8720
rect 2378 8686 2536 8720
rect 2570 8686 2586 8720
rect 182 8578 198 8612
rect 232 8578 390 8612
rect 424 8578 582 8612
rect 616 8578 774 8612
rect 808 8578 966 8612
rect 1000 8578 1158 8612
rect 1192 8578 1208 8612
rect 1560 8578 1576 8612
rect 1610 8578 1768 8612
rect 1802 8578 1960 8612
rect 1994 8578 2152 8612
rect 2186 8578 2344 8612
rect 2378 8578 2536 8612
rect 2570 8578 2586 8612
rect 182 8068 296 8102
rect 330 8068 486 8102
rect 520 8068 678 8102
rect 712 8068 870 8102
rect 904 8068 1062 8102
rect 1096 8068 1208 8102
rect 1560 8068 1672 8102
rect 1706 8068 1864 8102
rect 1898 8068 2056 8102
rect 2090 8068 2248 8102
rect 2282 8068 2438 8102
rect 2472 8068 2586 8102
<< viali >>
rect 294 9196 328 9230
rect 486 9196 520 9230
rect 678 9196 712 9230
rect 870 9196 904 9230
rect 1062 9196 1096 9230
rect 1672 9196 1706 9230
rect 1864 9196 1898 9230
rect 2056 9196 2090 9230
rect 2248 9196 2282 9230
rect 2440 9196 2474 9230
rect 198 8686 232 8720
rect 390 8686 424 8720
rect 582 8686 616 8720
rect 774 8686 808 8720
rect 966 8686 1000 8720
rect 1158 8686 1192 8720
rect 1576 8686 1610 8720
rect 1768 8686 1802 8720
rect 1960 8686 1994 8720
rect 2152 8686 2186 8720
rect 2344 8686 2378 8720
rect 2536 8686 2570 8720
rect 198 8578 232 8612
rect 390 8578 424 8612
rect 582 8578 616 8612
rect 774 8578 808 8612
rect 966 8578 1000 8612
rect 1158 8578 1192 8612
rect 1576 8578 1610 8612
rect 1768 8578 1802 8612
rect 1960 8578 1994 8612
rect 2152 8578 2186 8612
rect 2344 8578 2378 8612
rect 2536 8578 2570 8612
rect 296 8068 330 8102
rect 486 8068 520 8102
rect 678 8068 712 8102
rect 870 8068 904 8102
rect 1062 8068 1096 8102
rect 1672 8068 1706 8102
rect 1864 8068 1898 8102
rect 2056 8068 2090 8102
rect 2248 8068 2282 8102
rect 2438 8068 2472 8102
<< metal1 >>
rect 182 9230 1208 9236
rect 182 9196 294 9230
rect 328 9196 486 9230
rect 520 9196 678 9230
rect 712 9196 870 9230
rect 904 9196 1062 9230
rect 1096 9196 1208 9230
rect 182 9190 1208 9196
rect 1560 9230 2586 9236
rect 1560 9196 1672 9230
rect 1706 9196 1864 9230
rect 1898 9196 2056 9230
rect 2090 9196 2248 9230
rect 2282 9196 2440 9230
rect 2474 9196 2586 9230
rect 1560 9190 2586 9196
rect 130 8998 140 9158
rect 194 8998 204 9158
rect 322 8998 332 9158
rect 386 8998 396 9158
rect 514 8998 524 9158
rect 578 8998 588 9158
rect 706 8998 716 9158
rect 770 8998 780 9158
rect 898 8998 908 9158
rect 962 8998 972 9158
rect 1090 8998 1100 9158
rect 1154 8998 1164 9158
rect 1604 8998 1614 9158
rect 1668 8998 1678 9158
rect 1796 8998 1806 9158
rect 1860 8998 1870 9158
rect 1988 8998 1998 9158
rect 2052 8998 2062 9158
rect 2180 8998 2190 9158
rect 2244 8998 2254 9158
rect 2372 8998 2382 9158
rect 2436 8998 2446 9158
rect 2564 8998 2574 9158
rect 2628 8998 2638 9158
rect 226 8758 236 8918
rect 290 8758 300 8918
rect 418 8758 428 8918
rect 482 8758 492 8918
rect 610 8758 620 8918
rect 674 8758 684 8918
rect 802 8758 812 8918
rect 866 8758 876 8918
rect 994 8758 1004 8918
rect 1058 8758 1068 8918
rect 1186 8758 1196 8918
rect 1250 8758 1260 8918
rect 1508 8758 1518 8918
rect 1572 8758 1582 8918
rect 1700 8758 1710 8918
rect 1764 8758 1774 8918
rect 1892 8758 1902 8918
rect 1956 8758 1966 8918
rect 2084 8758 2094 8918
rect 2148 8758 2158 8918
rect 2276 8758 2286 8918
rect 2340 8758 2350 8918
rect 2468 8758 2478 8918
rect 2532 8758 2542 8918
rect 182 8720 1208 8726
rect 182 8686 198 8720
rect 232 8686 390 8720
rect 424 8686 582 8720
rect 616 8686 774 8720
rect 808 8686 966 8720
rect 1000 8686 1158 8720
rect 1192 8686 1208 8720
rect 182 8680 1208 8686
rect 1560 8720 2586 8726
rect 1560 8686 1576 8720
rect 1610 8686 1768 8720
rect 1802 8686 1960 8720
rect 1994 8686 2152 8720
rect 2186 8686 2344 8720
rect 2378 8686 2536 8720
rect 2570 8686 2586 8720
rect 1560 8680 2586 8686
rect 182 8612 1208 8618
rect 182 8578 198 8612
rect 232 8578 390 8612
rect 424 8578 582 8612
rect 616 8578 774 8612
rect 808 8578 966 8612
rect 1000 8578 1158 8612
rect 1192 8578 1208 8612
rect 182 8572 1208 8578
rect 1560 8612 2586 8618
rect 1560 8578 1576 8612
rect 1610 8578 1768 8612
rect 1802 8578 1960 8612
rect 1994 8578 2152 8612
rect 2186 8578 2344 8612
rect 2378 8578 2536 8612
rect 2570 8578 2586 8612
rect 1560 8572 2586 8578
rect 226 8380 236 8540
rect 290 8380 300 8540
rect 418 8380 428 8540
rect 482 8380 492 8540
rect 610 8380 620 8540
rect 674 8380 684 8540
rect 802 8380 812 8540
rect 866 8380 876 8540
rect 994 8380 1004 8540
rect 1058 8380 1068 8540
rect 1186 8380 1196 8540
rect 1250 8380 1260 8540
rect 1508 8380 1518 8540
rect 1572 8380 1582 8540
rect 1700 8380 1710 8540
rect 1764 8380 1774 8540
rect 1892 8380 1902 8540
rect 1956 8380 1966 8540
rect 2084 8380 2094 8540
rect 2148 8380 2158 8540
rect 2276 8380 2286 8540
rect 2340 8380 2350 8540
rect 2468 8380 2478 8540
rect 2532 8380 2542 8540
rect 130 8140 140 8300
rect 194 8140 204 8300
rect 322 8140 332 8300
rect 386 8140 396 8300
rect 514 8140 524 8300
rect 578 8140 588 8300
rect 706 8140 716 8300
rect 770 8140 780 8300
rect 898 8140 908 8300
rect 962 8140 972 8300
rect 1090 8140 1100 8300
rect 1154 8140 1164 8300
rect 1604 8140 1614 8300
rect 1668 8140 1678 8300
rect 1796 8140 1806 8300
rect 1860 8140 1870 8300
rect 1988 8140 1998 8300
rect 2052 8140 2062 8300
rect 2180 8140 2190 8300
rect 2244 8140 2254 8300
rect 2372 8140 2382 8300
rect 2436 8140 2446 8300
rect 2564 8140 2574 8300
rect 2628 8140 2638 8300
rect 182 8102 1208 8108
rect 182 8068 296 8102
rect 330 8068 486 8102
rect 520 8068 678 8102
rect 712 8068 870 8102
rect 904 8068 1062 8102
rect 1096 8068 1208 8102
rect 182 8062 1208 8068
rect 1560 8102 2586 8108
rect 1560 8068 1672 8102
rect 1706 8068 1864 8102
rect 1898 8068 2056 8102
rect 2090 8068 2248 8102
rect 2282 8068 2438 8102
rect 2472 8068 2586 8102
rect 1560 8062 2586 8068
<< via1 >>
rect 140 8998 194 9158
rect 332 8998 386 9158
rect 524 8998 578 9158
rect 716 8998 770 9158
rect 908 8998 962 9158
rect 1100 8998 1154 9158
rect 1614 8998 1668 9158
rect 1806 8998 1860 9158
rect 1998 8998 2052 9158
rect 2190 8998 2244 9158
rect 2382 8998 2436 9158
rect 2574 8998 2628 9158
rect 236 8758 290 8918
rect 428 8758 482 8918
rect 620 8758 674 8918
rect 812 8758 866 8918
rect 1004 8758 1058 8918
rect 1196 8758 1250 8918
rect 1518 8758 1572 8918
rect 1710 8758 1764 8918
rect 1902 8758 1956 8918
rect 2094 8758 2148 8918
rect 2286 8758 2340 8918
rect 2478 8758 2532 8918
rect 236 8380 290 8540
rect 428 8380 482 8540
rect 620 8380 674 8540
rect 812 8380 866 8540
rect 1004 8380 1058 8540
rect 1196 8380 1250 8540
rect 1518 8380 1572 8540
rect 1710 8380 1764 8540
rect 1902 8380 1956 8540
rect 2094 8380 2148 8540
rect 2286 8380 2340 8540
rect 2478 8380 2532 8540
rect 140 8140 194 8300
rect 332 8140 386 8300
rect 524 8140 578 8300
rect 716 8140 770 8300
rect 908 8140 962 8300
rect 1100 8140 1154 8300
rect 1614 8140 1668 8300
rect 1806 8140 1860 8300
rect 1998 8140 2052 8300
rect 2190 8140 2244 8300
rect 2382 8140 2436 8300
rect 2574 8140 2628 8300
<< metal2 >>
rect 140 9158 194 9168
rect 140 8988 194 8998
rect 332 9158 386 9168
rect 332 8988 386 8998
rect 524 9158 578 9168
rect 524 8988 578 8998
rect 716 9158 770 9168
rect 716 8988 770 8998
rect 908 9158 962 9168
rect 908 8988 962 8998
rect 1100 9158 1154 9168
rect 1100 8988 1154 8998
rect 1614 9158 1668 9168
rect 1614 8988 1668 8998
rect 1806 9158 1860 9168
rect 1806 8988 1860 8998
rect 1998 9158 2052 9168
rect 1998 8988 2052 8998
rect 2190 9158 2244 9168
rect 2190 8988 2244 8998
rect 2382 9158 2436 9168
rect 2382 8988 2436 8998
rect 2574 9158 2628 9168
rect 2574 8988 2628 8998
rect 236 8918 290 8928
rect 236 8748 290 8758
rect 428 8918 482 8928
rect 428 8748 482 8758
rect 620 8918 674 8928
rect 620 8748 674 8758
rect 812 8918 866 8928
rect 812 8748 866 8758
rect 1004 8918 1058 8928
rect 1004 8748 1058 8758
rect 1196 8918 1250 8928
rect 1196 8748 1250 8758
rect 1518 8918 1572 8928
rect 1518 8748 1572 8758
rect 1710 8918 1764 8928
rect 1710 8748 1764 8758
rect 1902 8918 1956 8928
rect 1902 8748 1956 8758
rect 2094 8918 2148 8928
rect 2094 8748 2148 8758
rect 2286 8918 2340 8928
rect 2286 8748 2340 8758
rect 2478 8918 2532 8928
rect 2478 8748 2532 8758
rect 236 8540 290 8550
rect 236 8370 290 8380
rect 428 8540 482 8550
rect 428 8370 482 8380
rect 620 8540 674 8550
rect 620 8370 674 8380
rect 812 8540 866 8550
rect 812 8370 866 8380
rect 1004 8540 1058 8550
rect 1004 8370 1058 8380
rect 1196 8540 1250 8550
rect 1196 8370 1250 8380
rect 1518 8540 1572 8550
rect 1518 8370 1572 8380
rect 1710 8540 1764 8550
rect 1710 8370 1764 8380
rect 1902 8540 1956 8550
rect 1902 8370 1956 8380
rect 2094 8540 2148 8550
rect 2094 8370 2148 8380
rect 2286 8540 2340 8550
rect 2286 8370 2340 8380
rect 2478 8540 2532 8550
rect 2478 8370 2532 8380
rect 140 8300 194 8310
rect 140 8130 194 8140
rect 332 8300 386 8310
rect 332 8130 386 8140
rect 524 8300 578 8310
rect 524 8130 578 8140
rect 716 8300 770 8310
rect 716 8130 770 8140
rect 908 8300 962 8310
rect 908 8130 962 8140
rect 1100 8300 1154 8310
rect 1100 8130 1154 8140
rect 1614 8300 1668 8310
rect 1614 8130 1668 8140
rect 1806 8300 1860 8310
rect 1806 8130 1860 8140
rect 1998 8300 2052 8310
rect 1998 8130 2052 8140
rect 2190 8300 2244 8310
rect 2190 8130 2244 8140
rect 2382 8300 2436 8310
rect 2382 8130 2436 8140
rect 2574 8300 2628 8310
rect 2574 8130 2628 8140
use sky130_fd_pr__nfet_01v8_lvt_324MKY  sky130_fd_pr__nfet_01v8_lvt_324MKY_0
timestamp 1647254192
transform 1 0 695 0 1 8649
box -695 -719 695 719
use sky130_fd_pr__nfet_01v8_lvt_324MKY  sky130_fd_pr__nfet_01v8_lvt_324MKY_2
timestamp 1647254192
transform -1 0 2073 0 1 8649
box -695 -719 695 719
<< end >>
