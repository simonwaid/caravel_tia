magic
tech sky130A
magscale 1 2
timestamp 1646993950
<< psubdiff >>
rect 8476 13900 8500 15280
rect 10040 13900 10064 15280
<< psubdiffcont >>
rect 8500 13900 10040 15280
<< locali >>
rect 8484 14040 8500 15280
rect -40 14020 8500 14040
rect -280 13900 8500 14020
rect 10040 14620 10056 15280
rect 10040 13900 11080 14620
rect -280 13760 11080 13900
rect 12442 13858 12652 13938
rect 12296 13760 12652 13858
rect -280 13460 12652 13760
rect -280 -2300 80 13460
rect 9900 13448 12652 13460
rect 9900 13440 12534 13448
rect 11060 13420 12440 13440
rect 12920 13380 13200 13440
rect 12900 8480 13220 13380
rect 18900 9790 19320 9800
rect 18900 9700 21010 9790
rect 12920 7330 13200 8480
rect 18900 7440 21010 7530
rect 12920 7320 13250 7330
rect 12920 7220 13340 7320
rect 12930 6180 13340 7220
rect 12930 6170 13260 6180
rect 12980 5000 13260 6170
rect 18880 5290 18930 5340
rect 18880 5200 20360 5290
rect 12910 4810 13280 5000
rect 12940 1720 13280 4810
rect 12910 1540 13280 1720
rect 18880 3010 18930 5200
rect 18880 2920 20360 3010
rect 12910 1340 18620 1540
rect 12880 1310 18620 1340
rect 12880 -860 13440 1310
rect 16580 -840 16820 1310
rect 18020 -1180 18620 1310
rect 13060 -2140 13220 -1360
rect 18260 -2140 18420 -1360
rect 18530 -1560 18620 -1180
rect 18880 760 18930 2920
rect 18880 670 20360 760
rect 18880 -1560 18930 670
rect -280 -2540 18540 -2300
rect 40 -2560 18540 -2540
rect 20760 -4780 21220 -4120
<< viali >>
rect 9300 13900 9800 15280
rect 17920 6300 18040 6480
rect 16446 5046 16624 5142
<< metal1 >>
rect 17670 15580 17680 15780
rect 17790 15580 17800 15780
rect 9294 15280 9806 15292
rect 9290 13900 9300 15280
rect 9800 13900 9810 15280
rect 12990 14600 13000 14720
rect 13080 14600 13090 14720
rect 17420 14360 17840 14480
rect 18000 14360 18010 14480
rect 12970 14080 12980 14200
rect 13060 14080 13070 14200
rect 13970 13980 13980 14100
rect 14100 14098 14140 14100
rect 14200 14098 14360 14100
rect 14100 13980 14360 14098
rect 14132 13976 14228 13980
rect 9294 13888 9806 13900
rect 12320 13740 12400 13800
rect 12320 13620 12520 13740
rect 12620 13620 12630 13740
rect 14900 11260 15040 13440
rect 17670 12400 17680 12580
rect 17980 12400 17990 12580
rect 17680 11480 17980 12400
rect 18800 11840 19020 11920
rect 18800 10980 18960 11840
rect 17420 10230 17540 10360
rect 14030 9840 14040 9980
rect 14180 9840 14360 9980
rect 18800 9920 18980 10980
rect 18800 9840 19040 9920
rect 18800 9660 18980 9840
rect 18800 9580 19040 9660
rect 18610 8500 18620 8760
rect 18800 7660 18980 9580
rect 12930 7180 13390 7240
rect 13430 7200 13610 7480
rect 17610 7400 17620 7660
rect 17800 7400 17810 7660
rect 18800 7580 19000 7660
rect 17620 7100 17800 7400
rect 18800 7310 18980 7580
rect 17914 6480 18046 6492
rect 12920 6250 13380 6310
rect 17910 6300 17920 6480
rect 18040 6300 18050 6480
rect 17914 6288 18046 6300
rect 16434 5142 16636 5148
rect 16434 5046 16446 5142
rect 16624 5046 16636 5142
rect 16434 5040 16636 5046
rect 14040 1340 14340 1800
rect 18210 1620 18220 2100
rect 18540 1620 18550 2100
rect 14040 -1310 14330 1340
rect 16290 580 16760 810
rect 18800 620 18980 5090
rect 18800 520 19020 620
rect 18800 490 18980 520
rect 14554 -4160 15600 -3240
rect 16420 -4160 16430 -3240
<< via1 >>
rect 17680 15580 17790 15780
rect 9300 13900 9800 15280
rect 13000 14600 13080 14720
rect 17840 14360 18000 14480
rect 12980 14080 13060 14200
rect 13980 13980 14100 14100
rect 12520 13620 12620 13740
rect 17680 12400 17980 12580
rect 14040 9840 14180 9980
rect 18620 8500 18800 8760
rect 17620 7400 17800 7660
rect 17920 6300 18040 6480
rect 16446 5046 16624 5142
rect 18220 1620 18540 2100
rect 15600 -4160 16420 -3240
<< metal2 >>
rect 17680 15780 17790 15790
rect 13060 15580 17680 15780
rect 17790 15580 21200 15780
rect 9300 15280 9800 15290
rect 13060 14730 13320 15580
rect 17680 15570 17790 15580
rect 18880 15560 19080 15580
rect 13000 14720 13320 14730
rect 13080 14600 13320 14720
rect 13760 15040 13880 15050
rect 13000 14590 13080 14600
rect 12980 14200 13060 14210
rect 13760 14200 13880 14900
rect 20920 15000 21200 15580
rect 18500 14520 18680 14536
rect 17640 14480 19080 14520
rect 17640 14360 17840 14480
rect 18000 14360 19080 14480
rect 17640 14320 19080 14360
rect 9800 13940 11260 14140
rect 13060 14080 13880 14200
rect 13980 14160 14520 14300
rect 13980 14100 14100 14160
rect 12980 14070 13060 14080
rect 9300 13890 9800 13900
rect 13980 13932 14100 13980
rect 13980 13790 14102 13932
rect 12520 13740 12620 13750
rect 13980 13720 14100 13790
rect 12520 13610 12620 13620
rect 13040 13500 14100 13720
rect 13040 9480 13720 13500
rect 17680 12580 17980 12590
rect 17680 12390 17980 12400
rect 13260 9240 13720 9480
rect 13860 11140 14060 11150
rect 14060 10900 14234 11140
rect 13860 10180 14234 10900
rect 18880 10560 19080 14320
rect 20920 12950 21180 15000
rect 20800 12940 21300 12950
rect 20800 12220 21300 12500
rect 20920 11600 21180 12220
rect 13860 10020 14380 10180
rect 13860 9980 14234 10020
rect 13860 9840 14040 9980
rect 14180 9840 14234 9980
rect 13040 9230 13260 9240
rect 13860 8306 14234 9840
rect 16800 8760 17020 8770
rect 17660 8760 18000 10380
rect 18620 8760 18800 8770
rect 18880 8760 19080 8940
rect 17020 8500 18620 8760
rect 18800 8500 19080 8760
rect 16800 8490 17020 8500
rect 17660 8480 18000 8500
rect 18620 8490 18800 8500
rect 13860 8120 14320 8306
rect 18880 8300 19080 8500
rect 12140 7760 12340 7770
rect 13220 7760 14320 8120
rect 12340 7560 12720 7760
rect 13140 7560 14320 7760
rect 20920 7780 21140 11600
rect 17620 7660 17800 7670
rect 12140 7550 12340 7560
rect 18240 7400 18520 7660
rect 17620 7390 17800 7400
rect 20920 7320 23100 7560
rect 12720 6920 13360 7120
rect 18360 7080 18680 7090
rect 18180 6800 18360 7080
rect 18180 6790 18680 6800
rect 17920 6480 18040 6490
rect 18180 6480 18660 6790
rect 17720 6300 17920 6480
rect 18040 6300 18660 6480
rect 17920 6290 18040 6300
rect 15840 5760 16380 6100
rect 16200 5140 16380 5760
rect 16446 5142 16624 5152
rect 16200 5046 16446 5140
rect 16200 5036 16624 5046
rect 16200 5020 16620 5036
rect 18220 2100 18540 2110
rect 18220 1610 18540 1620
rect 19160 1520 19300 6680
rect 22900 700 23100 7320
rect 20800 540 23100 700
rect 18040 160 18200 170
rect 18040 -50 18200 -40
rect 20800 -1360 21040 540
rect 16950 -1640 17820 -1400
rect 15600 -3240 16420 -3230
rect 15600 -4170 16420 -4160
rect 20760 -4240 21060 -4230
rect 20760 -4670 21060 -4660
<< via2 >>
rect 9300 13900 9800 15280
rect 13760 14900 13880 15040
rect 12520 13620 12620 13740
rect 17680 12400 17980 12580
rect 13040 9240 13260 9480
rect 13860 10900 14060 11140
rect 20800 12500 21300 12940
rect 16800 8500 17020 8760
rect 12140 7560 12340 7760
rect 20920 7560 21140 7780
rect 18360 6800 18680 7080
rect 18220 1620 18540 2100
rect 18040 -40 18200 160
rect 15600 -4160 16420 -3240
rect 20760 -4660 21060 -4240
<< metal3 >>
rect 9290 15280 9810 15285
rect 9290 13900 9300 15280
rect 9800 13900 9810 15280
rect 13750 15040 13890 15045
rect 13750 14900 13760 15040
rect 13880 14900 17000 15040
rect 13750 14895 13890 14900
rect 9290 13895 9810 13900
rect 12510 13740 12630 13745
rect 12510 13620 12520 13740
rect 12620 13620 14100 13740
rect 12510 13615 12630 13620
rect 12818 13500 14100 13620
rect 11850 11840 11860 11940
rect 12060 11840 12070 11940
rect 11380 7260 11680 7440
rect 9000 5840 9780 5980
rect 9000 4580 9860 5840
rect 9000 4420 9780 4580
rect 11870 1540 11880 11840
rect 12040 1540 12050 11840
rect 13860 11145 14060 13500
rect 13850 11140 14070 11145
rect 13850 10900 13860 11140
rect 14060 10900 14070 11140
rect 13850 10895 14070 10900
rect 13030 9480 13270 9485
rect 12480 9250 13040 9480
rect 12680 9240 13040 9250
rect 13260 9240 13270 9480
rect 13030 9235 13270 9240
rect 16820 8765 17000 14900
rect 20790 12940 21310 12945
rect 17840 12760 20800 12940
rect 17840 12585 17980 12760
rect 20790 12640 20800 12760
rect 17670 12580 17990 12585
rect 17670 12400 17680 12580
rect 17980 12568 17990 12580
rect 17980 12400 18000 12568
rect 20780 12500 20800 12640
rect 21300 12500 21310 12940
rect 17670 12395 17990 12400
rect 18880 11840 19080 12500
rect 20780 12495 21310 12500
rect 20780 12400 20980 12495
rect 16790 8760 17030 8765
rect 16790 8500 16800 8760
rect 17020 8500 17520 8760
rect 16790 8495 17030 8500
rect 20910 7780 21150 7785
rect 12130 7760 12350 7765
rect 12130 7560 12140 7760
rect 12340 7560 12350 7760
rect 12130 7555 12350 7560
rect 20910 7560 20920 7780
rect 21140 7560 21150 7780
rect 20910 7555 21150 7560
rect 18350 7080 18690 7085
rect 18350 6800 18360 7080
rect 18680 6800 18690 7080
rect 18350 6795 18690 6800
rect 18210 2100 18550 2105
rect 18210 1620 18220 2100
rect 18540 1620 18550 2100
rect 18210 1615 18550 1620
rect 18030 160 18210 165
rect 14900 -40 18040 160
rect 18200 -40 18210 160
rect 4100 -1730 9800 -700
rect 14900 -4000 15080 -40
rect 18030 -45 18210 -40
rect 15590 -3240 16430 -3235
rect 14554 -4800 15200 -4000
rect 15590 -4160 15600 -3240
rect 16420 -4160 16430 -3240
rect 15590 -4165 16430 -4160
rect 20750 -4240 21070 -4235
rect 20750 -4660 20760 -4240
rect 21060 -4660 21070 -4240
rect 20750 -4665 21070 -4660
<< via3 >>
rect 9300 13900 9800 15280
rect 11860 11840 12060 11940
rect 11880 1540 12040 11840
rect 20800 12500 21300 12940
rect 20920 7560 21140 7780
rect 18220 1620 18540 2100
rect 15600 -4160 16420 -3240
rect 20760 -4660 21060 -4240
<< metal4 >>
rect 9299 15280 9801 15281
rect 9299 13900 9300 15280
rect 9800 13900 9801 15280
rect 9299 13899 9801 13900
rect 20799 12940 21301 12941
rect 20799 12500 20800 12940
rect 21300 12500 21301 12940
rect 20799 12499 21301 12500
rect 20800 12380 21300 12499
rect 11859 11940 12061 11941
rect 11859 11840 11860 11940
rect 12060 11840 12061 11940
rect 11859 11839 11880 11840
rect 11879 8300 11880 11839
rect 12040 11839 12061 11840
rect 12040 8300 12041 11839
rect 20800 11820 21300 12220
rect 20900 7780 21400 8280
rect 9000 5840 9780 5980
rect 11879 5900 11880 7600
rect 12040 5900 12041 7600
rect 20900 7560 20920 7780
rect 21140 7560 21400 7780
rect 20900 7320 21400 7560
rect 9000 4800 9860 5840
rect 11879 1540 11880 5200
rect 12040 1540 12041 5200
rect 18219 2100 18541 2101
rect 18219 1620 18220 2100
rect 18540 1620 18541 2100
rect 18219 1619 18541 1620
rect 11879 1539 12041 1540
rect 11900 -1374 13900 -1300
rect 15599 -3240 16421 -3239
rect 15599 -4160 15600 -3240
rect 16420 -4160 16421 -3240
rect 15599 -4161 16421 -4160
rect 20759 -4240 21061 -4239
rect 20759 -4660 20760 -4240
rect 21060 -4660 21061 -4240
rect 20759 -4661 21061 -4660
<< via4 >>
rect 9300 13900 9800 15280
rect 20800 12500 21300 12940
rect 11720 7600 11880 8300
rect 11880 7600 12040 8300
rect 12040 7600 12320 8300
rect 11700 5200 11880 5900
rect 11880 5200 12040 5900
rect 12040 5200 12300 5900
rect 18220 1620 18540 2100
rect 15600 -4160 16420 -3240
rect 20760 -4660 21060 -4240
<< metal5 >>
rect 9276 15280 9824 15304
rect 9276 13900 9300 15280
rect 9800 13900 9824 15280
rect 9276 13876 9824 13900
rect 9300 12700 9800 13876
rect 20776 12940 21324 12964
rect 9300 12300 12900 12700
rect 20776 12500 20800 12940
rect 21300 12500 21324 12940
rect 20776 12476 21324 12500
rect 9300 11200 9800 12300
rect 10260 7200 10920 11780
rect 11700 8324 12300 12300
rect 11696 8300 12344 8324
rect 11696 7600 11720 8300
rect 12320 7600 12344 8300
rect 11696 7576 12344 7600
rect 20800 7320 21300 12476
rect 20800 7200 21400 7320
rect 10260 6300 21400 7200
rect 9000 5840 9780 5980
rect 9000 4580 9860 5840
rect 9000 4420 9780 4580
rect 8600 -2800 9800 -700
rect 10260 -1300 10920 6300
rect 11676 5900 12324 5924
rect 11676 5200 11700 5900
rect 12300 5200 12324 5900
rect 11676 5176 12324 5200
rect 11700 100 12300 5176
rect 18000 2100 18700 2300
rect 18000 1620 18220 2100
rect 18540 1620 18700 2100
rect 18000 100 18700 1620
rect 11700 -700 18700 100
rect 10260 -2240 17620 -1300
rect 11876 -2324 13924 -2240
rect 8600 -3216 16400 -2800
rect 8600 -3240 16444 -3216
rect 8600 -4160 15600 -3240
rect 16420 -4160 16444 -3240
rect 8600 -4184 16444 -4160
rect 8600 -4200 16400 -4184
rect 15600 -4800 16400 -4200
rect 16800 -4800 17600 -2240
rect 18000 -2900 18700 -700
rect 18000 -3600 21080 -2900
rect 20680 -4216 21080 -3600
rect 20680 -4240 21084 -4216
rect 20680 -4660 20760 -4240
rect 21060 -4660 21084 -4240
rect 20680 -4680 21084 -4660
rect 20736 -4684 21084 -4680
use isource_cmirror#0  isource_cmirror_2
timestamp 1646743514
transform 1 0 18900 0 1 9740
box 0 0 2044 2280
use isource_cmirror#0  isource_cmirror_3
timestamp 1646743514
transform 1 0 18900 0 1 7480
box 0 0 2044 2280
use isource_conv  isource_conv_0
timestamp 1646921651
transform 1 0 9200 0 1 -6200
box 3980 6900 13920 13860
use isource_conv_tsmal_nwell  isource_conv_tsmal_nwell_0
timestamp 1646921651
transform 1 0 12044 0 1 -1430
box 4070 6210 5960 9050
use isource_diffamp  isource_diffamp_0
timestamp 1646921651
transform 1 0 -280 0 1 16996
box 14560 -8200 18240 -5200
use isource_diffamp  isource_diffamp_1
timestamp 1646921651
transform 1 0 -280 0 1 21120
box 14560 -8200 18240 -5200
use isource_out  isource_out_0
timestamp 1646993950
transform 1 0 -4300 0 1 -13810
box 4320 8980 25514 15188
use isource_ref  isource_ref_0
timestamp 1646921651
transform 1 0 20 0 1 40
box -30 -40 13220 13420
use isource_startup  isource_startup_0
timestamp 1646921651
transform 1 0 10820 0 1 13700
box 200 0 2352 1238
use sky130_fd_pr__cap_mim_m3_1_WXTTNJ#0  sky130_fd_pr__cap_mim_m3_1_WXTTNJ_0
timestamp 1646921651
transform 1 0 19490 0 1 10040
box -2150 -2100 2149 2100
use sky130_fd_pr__cap_mim_m3_2_LJ5JLG#1  sky130_fd_pr__cap_mim_m3_2_LJ5JLG_0
timestamp 1646921651
transform 1 0 7151 0 1 1700
box -3351 -3101 3373 3101
use sky130_fd_pr__cap_mim_m3_2_LJ5JLG#1  sky130_fd_pr__cap_mim_m3_2_LJ5JLG_1
timestamp 1646921651
transform 1 0 7151 0 1 8700
box -3351 -3101 3373 3101
<< labels >>
rlabel metal3 14600 -4600 15000 -4200 7 I_ref
port 2 w
rlabel metal1 14040 730 14330 920 1 VM3G
rlabel metal2 17660 -1630 17810 -1400 3 VM3D
rlabel metal1 16290 580 16490 800 3 VM22D
rlabel metal3 11380 7260 11680 7440 1 VM12D
rlabel metal1 13440 7380 13580 7460 1 VM12G
rlabel metal5 16940 -4640 17440 -4120 1 VP
port 1 n
rlabel metal5 15800 -4600 16200 -4200 1 VN
port 3 n
rlabel metal2 13720 7620 14040 8060 1 VM11D
rlabel metal2 18260 7400 18480 7660 1 VM14D
rlabel metal1 14908 12062 15034 12202 1 VM9D
rlabel metal2 17100 8540 17460 8740 1 VM8D
rlabel metal2 13280 12860 13440 13080 1 VM2D
<< end >>
