magic
tech sky130A
magscale 1 2
timestamp 1647254192
<< locali >>
rect 40 4820 12900 4940
rect 20 3600 12880 3720
rect 40 2380 12900 2500
rect 40 1160 12900 1280
<< viali >>
rect 20 1440 80 1640
rect 12820 1440 12900 1640
<< metal1 >>
rect 12450 4720 12460 4800
rect 12660 4720 12670 4800
rect 12450 3740 12460 3820
rect 12660 3740 12670 3820
rect 12450 3480 12460 3560
rect 12660 3480 12670 3560
rect 12450 2520 12460 2600
rect 12660 2520 12670 2600
rect 12450 2220 12460 2300
rect 12660 2220 12670 2300
rect 14 1640 86 1652
rect 12814 1640 12906 1652
rect 14 1440 20 1640
rect 80 1440 180 1640
rect 12720 1440 12820 1640
rect 12900 1440 12906 1640
rect 14 1428 86 1440
rect 12814 1428 12906 1440
rect 12450 1300 12460 1380
rect 12660 1300 12670 1380
rect 12450 1060 12460 1140
rect 12660 1060 12670 1140
rect 12470 80 12480 160
rect 12680 80 12690 160
<< via1 >>
rect 12460 4720 12660 4800
rect 12460 3740 12660 3820
rect 12460 3480 12660 3560
rect 12460 2520 12660 2600
rect 12460 2220 12660 2300
rect 12460 1300 12660 1380
rect 12460 1060 12660 1140
rect 12480 80 12680 160
<< metal2 >>
rect 12460 4800 12660 4810
rect 12460 4710 12660 4720
rect 12120 4580 12320 4590
rect 12120 4510 12320 4520
rect 220 4020 520 4030
rect 220 3950 520 3960
rect 12460 3820 12660 3830
rect 12460 3730 12660 3740
rect 12460 3560 12660 3570
rect 12460 3470 12660 3480
rect 12120 3360 12320 3370
rect 12120 3290 12320 3300
rect 220 2800 520 2810
rect 220 2730 520 2740
rect 12460 2600 12660 2610
rect 12460 2510 12660 2520
rect 12460 2300 12660 2310
rect 12460 2210 12660 2220
rect 12460 2140 12660 2150
rect 12460 2070 12660 2080
rect 620 1560 920 1570
rect 620 1490 920 1500
rect 12460 1380 12660 1390
rect 12460 1290 12660 1300
rect 12460 1140 12660 1150
rect 12460 1050 12660 1060
rect 12120 920 12320 930
rect 12120 850 12320 860
rect 220 340 520 350
rect 220 270 520 280
rect 12480 160 12680 170
rect 12480 70 12680 80
<< via2 >>
rect 12460 4720 12660 4800
rect 12120 4520 12320 4580
rect 220 3960 520 4020
rect 12460 3740 12660 3820
rect 12460 3480 12660 3560
rect 12120 3300 12320 3360
rect 220 2740 520 2800
rect 12460 2520 12660 2600
rect 12460 2220 12660 2300
rect 12460 2080 12660 2140
rect 620 1500 920 1560
rect 12460 1300 12660 1380
rect 12460 1060 12660 1140
rect 12120 860 12320 920
rect 220 280 520 340
rect 12480 80 12680 160
<< metal3 >>
rect 210 4020 530 4025
rect 210 3960 220 4020
rect 520 3960 530 4020
rect 210 3955 530 3960
rect 220 2805 520 3955
rect 210 2800 530 2805
rect 210 2740 220 2800
rect 520 2740 530 2800
rect 210 2735 530 2740
rect 220 345 520 2735
rect 620 1565 920 4940
rect 12460 4805 12660 4940
rect 12450 4800 12670 4805
rect 12450 4720 12460 4800
rect 12660 4720 12670 4800
rect 12450 4715 12670 4720
rect 12110 4580 12330 4585
rect 12110 4520 12120 4580
rect 12320 4520 12330 4580
rect 12110 4515 12330 4520
rect 12120 3365 12320 4515
rect 12460 3825 12660 4715
rect 12450 3820 12670 3825
rect 12450 3740 12460 3820
rect 12660 3740 12670 3820
rect 12450 3735 12670 3740
rect 12460 3565 12660 3735
rect 12450 3560 12670 3565
rect 12450 3480 12460 3560
rect 12660 3480 12670 3560
rect 12450 3475 12670 3480
rect 12110 3360 12330 3365
rect 12110 3300 12120 3360
rect 12320 3300 12330 3360
rect 12110 3295 12330 3300
rect 610 1560 930 1565
rect 610 1500 620 1560
rect 920 1500 930 1560
rect 610 1495 930 1500
rect 12120 925 12320 3295
rect 12460 2605 12660 3475
rect 12450 2600 12670 2605
rect 12450 2520 12460 2600
rect 12660 2520 12670 2600
rect 12450 2515 12670 2520
rect 12460 2305 12660 2515
rect 12450 2300 12670 2305
rect 12450 2220 12460 2300
rect 12660 2220 12670 2300
rect 12450 2215 12670 2220
rect 12460 2145 12660 2215
rect 12450 2140 12670 2145
rect 12450 2080 12460 2140
rect 12660 2080 12670 2140
rect 12450 2075 12670 2080
rect 12460 1385 12660 2075
rect 12450 1380 12670 1385
rect 12450 1300 12460 1380
rect 12660 1300 12670 1380
rect 12450 1295 12670 1300
rect 12460 1145 12660 1295
rect 12450 1140 12670 1145
rect 12450 1060 12460 1140
rect 12660 1060 12670 1140
rect 12450 1055 12670 1060
rect 12110 920 12330 925
rect 12110 860 12120 920
rect 12320 860 12330 920
rect 12110 855 12330 860
rect 210 340 530 345
rect 210 280 220 340
rect 520 280 530 340
rect 210 275 530 280
rect 12460 165 12660 1055
rect 12460 160 12690 165
rect 12460 80 12480 160
rect 12680 80 12690 160
rect 12460 75 12690 80
rect 12460 40 12660 75
use isource_ref_transistor  isource_ref_transistor_0
timestamp 1647254192
transform 1 0 493 0 1 117
box -493 -117 12421 1103
use isource_ref_transistor  isource_ref_transistor_1
timestamp 1647254192
transform 1 0 493 0 1 1337
box -493 -117 12421 1103
use isource_ref_transistor  isource_ref_transistor_3
timestamp 1647254192
transform 1 0 493 0 1 2557
box -493 -117 12421 1103
use isource_ref_transistor  isource_ref_transistor_4
timestamp 1647254192
transform 1 0 493 0 1 3777
box -493 -117 12421 1103
<< end >>
