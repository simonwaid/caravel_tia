* SPICE3 file created from isource.ext - technology: sky130A

.subckt isource I_ref VN VP
X0 VP VM8D sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X1 VM12G VM14D VP VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.75622e+14p ps=1.58256e+09u w=4e+06u l=150000u
X2 VM12G VM14D VP VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3 VP VM14D VM12G VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4 VM12G VM14D VP VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5 VP VM14D VM12G VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6 VM12G VM14D VP VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7 VM12G VM14D VP VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8 VP VM14D VM12G VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9 VP VM14D VM12G VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10 VP VM14D VM12G VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X11 VM12G VM14D VP VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X12 VM12G VM14D VP VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X13 VP VM14D VM12G VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X14 VM12G VM14D VP VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X15 VM12G VM14D VP VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X16 VP VM14D VM12G VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X17 VP VM14D VM12G VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X18 VP VM14D VM12G VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X19 VP VM14D VM12G VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X20 VM12G VM14D VP VM12G sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X21 VP VM11D isource_startup_0/m1_330_800# VP sky130_fd_pr__pfet_01v8 ad=6.18049e+13p pd=4.649e+08u as=0p ps=0u w=500000u l=2e+06u
X22 VM8D isource_startup_0/m1_330_800# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.4945e+13p ps=2.5898e+08u w=500000u l=2e+06u
X23 VN VM11D isource_startup_0/m1_330_800# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X24 isource_startup_0/m1_330_800# VM11D VN VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X25 isource_startup_0/m1_330_800# VM11D VN VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X26 VN VM11D isource_startup_0/m1_330_800# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X27 VN VM11D isource_startup_0/m1_330_800# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X28 isource_startup_0/m1_330_800# VM11D VN VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X29 isource_startup_0/m1_330_800# VM11D VN VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X30 isource_startup_0/m1_330_800# VM11D VN VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X31 VN VM11D isource_startup_0/m1_330_800# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X32 VN VM11D isource_startup_0/m1_330_800# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X33 VN VM2D VM2D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X34 VM2D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X35 VM2D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X36 VN VM2D VM2D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X37 VM2D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X38 VN VM2D VM2D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X39 VN VM2D VM2D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X40 VN VM2D VM2D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X41 VM2D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X42 VM2D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X43 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X44 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X45 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X46 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X47 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X48 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X49 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X50 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X51 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X52 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X53 VN VM2D VM2D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X54 VM2D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X55 VM2D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X56 VN VM2D VM2D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X57 VM2D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X58 VN VM2D VM2D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X59 VN VM2D VM2D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X60 VN VM2D VM2D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X61 VM2D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X62 VM2D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X63 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X64 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X65 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X66 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X67 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X68 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X69 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X70 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X71 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X72 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X73 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X74 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X75 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X76 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X77 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X78 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X79 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X80 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X81 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X82 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X83 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X84 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X85 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X86 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X87 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X88 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X89 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X90 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X91 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X92 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X93 VN VM2D VM2D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X94 VM2D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X95 VM2D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X96 VN VM2D VM2D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X97 VM2D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X98 VN VM2D VM2D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X99 VN VM2D VM2D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X100 VN VM2D VM2D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X101 VM2D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X102 VM2D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X103 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X104 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X105 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X106 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X107 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X108 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X109 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X110 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X111 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X112 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X113 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X114 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X115 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X116 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X117 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X118 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X119 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X120 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X121 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X122 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X123 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X124 VM12D VM2D VM11D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X125 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X126 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X127 VM11D VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X128 VM12D VM12G VN isource_ref_0/sky130_fd_pr__nfet_01v8_WY4VMC_0/a_n1389_n574# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X129 VN VM12G VM12D isource_ref_0/sky130_fd_pr__nfet_01v8_WY4VMC_0/a_n1389_n574# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X130 isource_cmirror_2/m1_250_820# VM8D VM9D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X131 isource_cmirror_2/m1_250_820# VM8D VM9D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X132 VP VM8D isource_cmirror_2/m1_250_820# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X133 VP VM8D isource_cmirror_2/m1_250_820# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X134 isource_cmirror_2/m1_250_820# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X135 VP VM8D isource_cmirror_2/m1_250_820# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X136 VP VM8D isource_cmirror_2/m1_250_820# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X137 isource_cmirror_2/m1_250_820# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X138 VP VM8D isource_cmirror_2/m1_250_820# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X139 VP VM8D isource_cmirror_2/m1_250_820# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X140 isource_cmirror_2/m1_250_820# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X141 isource_cmirror_2/m1_250_820# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X142 isource_cmirror_3/m1_250_820# VM8D VM8D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X143 isource_cmirror_3/m1_250_820# VM8D VM8D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X144 VP VM8D isource_cmirror_3/m1_250_820# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X145 VP VM8D isource_cmirror_3/m1_250_820# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X146 isource_cmirror_3/m1_250_820# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X147 VP VM8D isource_cmirror_3/m1_250_820# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X148 VP VM8D isource_cmirror_3/m1_250_820# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X149 isource_cmirror_3/m1_250_820# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X150 VP VM8D isource_cmirror_3/m1_250_820# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X151 VP VM8D isource_cmirror_3/m1_250_820# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X152 isource_cmirror_3/m1_250_820# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X153 isource_cmirror_3/m1_250_820# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X154 m2_19160_1520# VM8D VM14D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X155 m2_19160_1520# VM8D VM14D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X156 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X157 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X158 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X159 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X160 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X161 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X162 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X163 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X164 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X165 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X166 m2_19160_1520# VM8D VM14D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X167 m2_19160_1520# VM8D VM14D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X168 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X169 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X170 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X171 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X172 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X173 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X174 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X175 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X176 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X177 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X178 m2_19160_1520# VM8D VM14D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X179 m2_19160_1520# VM8D VM14D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X180 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X181 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X182 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X183 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X184 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X185 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X186 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X187 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X188 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X189 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X190 m2_19160_1520# VM8D VM14D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X191 m2_19160_1520# VM8D VM14D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X192 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X193 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X194 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X195 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X196 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X197 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X198 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X199 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X200 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X201 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X202 m2_19160_1520# VM8D VM14D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X203 m2_19160_1520# VM8D VM14D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X204 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X205 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X206 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X207 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X208 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X209 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X210 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X211 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X212 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X213 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X214 m2_19160_1520# VM8D VM14D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X215 m2_19160_1520# VM8D VM14D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X216 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X217 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X218 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X219 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X220 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X221 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X222 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X223 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X224 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X225 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X226 isource_conv_0/m1_7960_7820# isource_conv_0/m1_7420_10260# VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X227 isource_conv_0/m1_6900_7820# isource_conv_0/m1_7420_10260# VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X228 VM3G isource_conv_0/m1_5300_10260# VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X229 isource_conv_0/m1_5840_7820# isource_conv_0/m1_5300_10260# VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X230 isource_conv_0/m1_5840_7820# isource_conv_0/m1_6360_10260# VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X231 VN isource_conv_0/m1_8480_10260# VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X232 isource_conv_0/m1_6900_7820# isource_conv_0/m1_6360_10260# VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X233 isource_conv_0/m1_7960_7820# isource_conv_0/m1_8480_10260# VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X234 VM14D VM12G VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X235 VN VM12G VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X236 VM3G isource_conv_0/m1_4160_10260# VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X237 VM12G isource_conv_0/m1_4160_10260# VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X238 VM11D VM9D VM8D VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X239 VM11D VM9D VM8D VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X240 VM8D VM9D VM11D VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X241 VM8D VM9D VM11D VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X242 VM11D VM9D VM8D VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X243 VM8D VM9D VM11D VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X244 VM11D VM9D VM8D VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X245 VM8D VM9D VM11D VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X246 VM11D VM9D VM8D VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X247 VM8D VM9D VM11D VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X248 VM11D VM9D VM8D VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X249 VM11D VM9D VM8D VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X250 VM8D VM9D VM11D VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X251 VM8D VM9D VM11D VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X252 VM8D VM9D VM11D VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X253 VM11D VM9D VM8D VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X254 VM11D VM9D VM8D VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X255 VM8D VM9D VM11D VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X256 VM11D VM9D VM8D VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X257 VM8D VM9D VM11D VM11D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X258 VM2D VM9D VM9D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X259 VM2D VM9D VM9D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X260 VM9D VM9D VM2D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X261 VM9D VM9D VM2D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X262 VM2D VM9D VM9D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X263 VM9D VM9D VM2D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X264 VM2D VM9D VM9D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X265 VM9D VM9D VM2D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X266 VM2D VM9D VM9D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X267 VM9D VM9D VM2D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X268 VM2D VM9D VM9D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X269 VM2D VM9D VM9D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X270 VM9D VM9D VM2D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X271 VM9D VM9D VM2D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X272 VM9D VM9D VM2D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X273 VM2D VM9D VM9D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X274 VM2D VM9D VM9D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X275 VM9D VM9D VM2D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X276 VM2D VM9D VM9D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X277 VM9D VM9D VM2D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X278 VN VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X279 VN VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X280 a_19136_n1351# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X281 I_ref VM22D a_216_n2258# VN sky130_fd_pr__nfet_01v8_lvt ad=1.552e+13p pd=1.0376e+08u as=0p ps=0u w=4e+06u l=150000u
X282 VM3D a_216_n2258# VM22D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X283 VP VM8D a_19136_n1351# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X284 a_18646_n4664# a_19176_n2232# VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X285 VM3D a_216_n2258# VM22D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X286 VM22D a_216_n2258# VM3D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X287 VM22D a_216_n2258# VM3D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X288 VM22D a_216_n2258# VM3D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X289 a_19136_n1351# VM8D VM22D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X290 VN a_20236_n2232# VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X291 VM3D a_216_n2258# VM22D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X292 I_ref VM22D a_216_n2258# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X293 VM3D a_216_n2258# VM22D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X294 a_19706_n4664# a_19176_n2232# VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X295 VM3D VM3G VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X296 a_216_n2258# VM22D I_ref VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X297 a_216_n2258# VM22D I_ref VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X298 VP VM8D a_19136_n1351# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X299 a_19706_n4664# a_20236_n2232# VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X300 I_ref VM22D a_216_n2258# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X301 a_18646_n4664# a_216_n2258# VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X302 I_ref VM22D a_216_n2258# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X303 a_216_n2258# VM22D I_ref VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X304 a_216_n2258# VM22D I_ref VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X305 I_ref VM22D a_216_n2258# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X306 I_ref VM22D a_216_n2258# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X307 VM3D VM3G VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X308 I_ref VM22D a_216_n2258# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X309 a_216_n2258# VM22D I_ref VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X310 a_216_n2258# VM22D I_ref VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X311 I_ref VM22D a_216_n2258# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X312 I_ref VM22D a_216_n2258# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X313 a_19136_n1351# VM8D VM22D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X314 a_19136_n1351# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X315 VN VM3G VM3D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X316 VM3D a_216_n2258# VM22D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X317 a_19136_n1351# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X318 VP VM8D a_19136_n1351# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X319 a_216_n2258# VM22D I_ref VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X320 VM22D a_216_n2258# VM3D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X321 VN VM3G VM3D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X322 I_ref VM22D a_216_n2258# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X323 a_216_n2258# VM22D I_ref VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X324 VP VM8D a_19136_n1351# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X325 VM3D a_216_n2258# VM22D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X326 VM3D a_216_n2258# VM22D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X327 VP VM8D a_19136_n1351# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X328 VM22D a_216_n2258# VM3D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X329 VM3D a_216_n2258# VM22D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X330 VM22D a_216_n2258# VM3D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X331 a_216_n2258# VM22D I_ref VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X332 VM3D a_216_n2258# VM22D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X333 VM22D a_216_n2258# VM3D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X334 VM22D a_216_n2258# VM3D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X335 VM22D a_216_n2258# VM3D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X336 a_19136_n1351# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X337 VM3D a_216_n2258# VM22D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X338 VM22D a_216_n2258# VM3D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X339 a_216_n2258# VM22D I_ref VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X340 VP VM8D a_19136_n1351# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
.ends
