* SPICE3 file created from esd-array.ext - technology: sky130A

D0 VSUBS m1_n9090_410# sky130_fd_pr__diode_pw2nd_05v5 pj=8e+06u area=4e+12p
D1 VSUBS m1_n9090_410# sky130_fd_pr__diode_pw2nd_05v5 pj=8e+06u area=4e+12p
D2 VSUBS m1_n9090_410# sky130_fd_pr__diode_pw2nd_05v5 pj=8e+06u area=4e+12p
D3 VSUBS m1_n9090_410# sky130_fd_pr__diode_pw2nd_05v5 pj=8e+06u area=4e+12p
D4 VSUBS m1_n9090_410# sky130_fd_pr__diode_pw2nd_05v5 pj=8e+06u area=4e+12p
D5 VSUBS m1_n9090_410# sky130_fd_pr__diode_pw2nd_05v5 pj=8e+06u area=4e+12p
D6 VSUBS m1_n9090_410# sky130_fd_pr__diode_pw2nd_05v5 pj=8e+06u area=4e+12p
D7 VSUBS m1_n9090_410# sky130_fd_pr__diode_pw2nd_05v5 pj=8e+06u area=4e+12p
D8 VSUBS m1_n9090_410# sky130_fd_pr__diode_pw2nd_05v5 pj=8e+06u area=4e+12p
D9 VSUBS m1_n9090_410# sky130_fd_pr__diode_pw2nd_05v5 pj=8e+06u area=4e+12p
D10 m1_n9090_410# w_n9230_1690# sky130_fd_pr__diode_pd2nw_05v5 pj=8e+06u area=4e+12p
D11 m1_n9090_410# w_n9230_1690# sky130_fd_pr__diode_pd2nw_05v5 pj=8e+06u area=4e+12p
D12 m1_n9090_410# w_n9230_1690# sky130_fd_pr__diode_pd2nw_05v5 pj=8e+06u area=4e+12p
D13 m1_n9090_410# w_n9230_1690# sky130_fd_pr__diode_pd2nw_05v5 pj=8e+06u area=4e+12p
D14 m1_n9090_410# w_n9230_1690# sky130_fd_pr__diode_pd2nw_05v5 pj=8e+06u area=4e+12p
D15 m1_n9090_410# w_n9230_1690# sky130_fd_pr__diode_pd2nw_05v5 pj=8e+06u area=4e+12p
D16 m1_n9090_410# w_n9230_1690# sky130_fd_pr__diode_pd2nw_05v5 pj=8e+06u area=4e+12p
D17 m1_n9090_410# w_n9230_1690# sky130_fd_pr__diode_pd2nw_05v5 pj=8e+06u area=4e+12p
D18 m1_n9090_410# w_n9230_1690# sky130_fd_pr__diode_pd2nw_05v5 pj=8e+06u area=4e+12p
D19 m1_n9090_410# w_n9230_1690# sky130_fd_pr__diode_pd2nw_05v5 pj=8e+06u area=4e+12p
