magic
tech sky130A
magscale 1 2
timestamp 1647254192
<< pwell >>
rect 10 5090 1860 5220
<< locali >>
rect 0 7770 1870 7840
rect 0 5220 70 7770
rect 1800 5220 1870 7770
rect 0 5210 1870 5220
rect 0 5140 1020 5210
rect 1730 5150 1870 5210
rect 1730 5140 2860 5150
rect 0 5080 2860 5140
rect 0 70 70 5080
rect 2790 70 2860 5080
rect 0 40 2860 70
rect 0 0 990 40
rect 980 -70 990 0
rect 1950 0 2860 40
rect 1950 -70 1960 0
<< viali >>
rect 1020 5140 1730 5210
rect 990 -70 1950 40
<< metal1 >>
rect 0 7660 1870 7750
rect 0 7190 100 7660
rect 130 7460 140 7620
rect 200 7460 210 7620
rect 320 7460 330 7620
rect 390 7460 400 7620
rect 510 7460 520 7620
rect 580 7460 590 7620
rect 700 7460 710 7620
rect 770 7460 780 7620
rect 900 7460 910 7620
rect 970 7460 980 7620
rect 1090 7460 1100 7620
rect 1160 7460 1170 7620
rect 1280 7460 1290 7620
rect 1350 7460 1360 7620
rect 1470 7460 1480 7620
rect 1540 7460 1550 7620
rect 1660 7460 1670 7620
rect 1730 7460 1740 7620
rect 220 7220 230 7380
rect 290 7220 300 7380
rect 420 7220 430 7380
rect 490 7220 500 7380
rect 610 7220 620 7380
rect 680 7220 690 7380
rect 800 7220 810 7380
rect 870 7220 880 7380
rect 990 7220 1000 7380
rect 1060 7220 1070 7380
rect 1180 7220 1190 7380
rect 1250 7220 1260 7380
rect 1380 7220 1390 7380
rect 1450 7220 1460 7380
rect 1570 7220 1580 7380
rect 1640 7220 1650 7380
rect 1770 7190 1870 7660
rect 0 7040 1870 7190
rect 0 6570 100 7040
rect 220 6850 230 7010
rect 290 6850 300 7010
rect 420 6850 430 7010
rect 490 6850 500 7010
rect 610 6850 620 7010
rect 680 6850 690 7010
rect 800 6850 810 7010
rect 870 6850 880 7010
rect 990 6850 1000 7010
rect 1060 6850 1070 7010
rect 1180 6850 1190 7010
rect 1250 6850 1260 7010
rect 1380 6850 1390 7010
rect 1450 6850 1460 7010
rect 1570 6850 1580 7010
rect 1640 6850 1650 7010
rect 130 6610 140 6770
rect 200 6610 210 6770
rect 320 6610 330 6770
rect 390 6610 400 6770
rect 510 6610 520 6770
rect 580 6610 590 6770
rect 700 6610 710 6770
rect 770 6610 780 6770
rect 900 6610 910 6770
rect 970 6610 980 6770
rect 1090 6610 1100 6770
rect 1160 6610 1170 6770
rect 1280 6610 1290 6770
rect 1350 6610 1360 6770
rect 1470 6610 1480 6770
rect 1540 6610 1550 6770
rect 1660 6610 1670 6770
rect 1730 6610 1740 6770
rect 1770 6570 1870 7040
rect 0 6420 1870 6570
rect 0 5960 100 6420
rect 130 6230 140 6390
rect 200 6230 210 6390
rect 320 6230 330 6390
rect 390 6230 400 6390
rect 510 6230 520 6390
rect 580 6230 590 6390
rect 700 6230 710 6390
rect 770 6230 780 6390
rect 900 6230 910 6390
rect 970 6230 980 6390
rect 1090 6230 1100 6390
rect 1160 6230 1170 6390
rect 1280 6230 1290 6390
rect 1350 6230 1360 6390
rect 1470 6230 1480 6390
rect 1540 6230 1550 6390
rect 1660 6230 1670 6390
rect 1730 6230 1740 6390
rect 220 5990 230 6150
rect 290 5990 300 6150
rect 420 5990 430 6150
rect 490 5990 500 6150
rect 610 5990 620 6150
rect 680 5990 690 6150
rect 800 5990 810 6150
rect 870 5990 880 6150
rect 990 5990 1000 6150
rect 1060 5990 1070 6150
rect 1180 5990 1190 6150
rect 1250 5990 1260 6150
rect 1380 5990 1390 6150
rect 1450 5990 1460 6150
rect 1570 5990 1580 6150
rect 1640 5990 1650 6150
rect 1770 5960 1870 6420
rect 0 5800 1870 5960
rect 0 5340 100 5800
rect 220 5610 230 5770
rect 290 5610 300 5770
rect 420 5610 430 5770
rect 490 5610 500 5770
rect 610 5610 620 5770
rect 680 5610 690 5770
rect 800 5610 810 5770
rect 870 5610 880 5770
rect 990 5610 1000 5770
rect 1060 5610 1070 5770
rect 1180 5610 1190 5770
rect 1250 5610 1260 5770
rect 1380 5610 1390 5770
rect 1450 5610 1460 5770
rect 1570 5610 1580 5770
rect 1640 5610 1650 5770
rect 130 5370 140 5530
rect 200 5370 210 5530
rect 320 5370 330 5530
rect 390 5370 400 5530
rect 510 5370 520 5530
rect 580 5370 590 5530
rect 700 5370 710 5530
rect 770 5370 780 5530
rect 900 5370 910 5530
rect 970 5370 980 5530
rect 1090 5370 1100 5530
rect 1160 5370 1170 5530
rect 1280 5370 1290 5530
rect 1350 5370 1360 5530
rect 1470 5370 1480 5530
rect 1540 5370 1550 5530
rect 1660 5370 1670 5530
rect 1730 5370 1740 5530
rect 1770 5340 1870 5800
rect 0 5250 1870 5340
rect 0 5090 100 5250
rect 1008 5210 1742 5216
rect 1008 5140 1020 5210
rect 1730 5140 1742 5210
rect 1008 5134 1742 5140
rect 1770 5090 1870 5250
rect 0 4970 2860 5090
rect 0 4500 100 4970
rect 130 4780 140 4940
rect 200 4780 210 4940
rect 440 4780 450 4940
rect 510 4780 520 4940
rect 760 4780 770 4940
rect 830 4780 840 4940
rect 1080 4780 1090 4940
rect 1150 4780 1160 4940
rect 1390 4780 1400 4940
rect 1460 4780 1470 4940
rect 1710 4780 1720 4940
rect 1780 4780 1790 4940
rect 2020 4780 2030 4940
rect 2090 4780 2100 4940
rect 2340 4780 2350 4940
rect 2410 4780 2420 4940
rect 2650 4780 2660 4940
rect 2720 4780 2730 4940
rect 280 4540 290 4700
rect 350 4540 360 4700
rect 600 4540 610 4700
rect 670 4540 680 4700
rect 920 4540 930 4700
rect 990 4540 1000 4700
rect 1230 4540 1240 4700
rect 1300 4540 1310 4700
rect 1550 4540 1560 4700
rect 1620 4540 1630 4700
rect 1860 4540 1870 4700
rect 1930 4540 1940 4700
rect 2180 4540 2190 4700
rect 2250 4540 2260 4700
rect 2500 4540 2510 4700
rect 2570 4540 2580 4700
rect 2760 4500 2860 4970
rect 0 4350 2860 4500
rect 0 3880 100 4350
rect 280 4160 290 4320
rect 350 4160 360 4320
rect 600 4160 610 4320
rect 670 4160 680 4320
rect 920 4160 930 4320
rect 990 4160 1000 4320
rect 1230 4160 1240 4320
rect 1300 4160 1310 4320
rect 1550 4160 1560 4320
rect 1620 4160 1630 4320
rect 1860 4160 1870 4320
rect 1930 4160 1940 4320
rect 2180 4160 2190 4320
rect 2250 4160 2260 4320
rect 2500 4160 2510 4320
rect 2570 4160 2580 4320
rect 130 3920 140 4080
rect 200 3920 210 4080
rect 440 3920 450 4080
rect 510 3920 520 4080
rect 760 3920 770 4080
rect 830 3920 840 4080
rect 1080 3920 1090 4080
rect 1150 3920 1160 4080
rect 1390 3920 1400 4080
rect 1460 3920 1470 4080
rect 1710 3920 1720 4080
rect 1780 3920 1790 4080
rect 2020 3920 2030 4080
rect 2090 3920 2100 4080
rect 2340 3920 2350 4080
rect 2410 3920 2420 4080
rect 2650 3920 2660 4080
rect 2720 3920 2730 4080
rect 2760 3880 2860 4350
rect 0 3730 2860 3880
rect 0 3260 100 3730
rect 130 3540 140 3700
rect 200 3540 210 3700
rect 440 3540 450 3700
rect 510 3540 520 3700
rect 760 3540 770 3700
rect 830 3540 840 3700
rect 1080 3540 1090 3700
rect 1150 3540 1160 3700
rect 1390 3540 1400 3700
rect 1460 3540 1470 3700
rect 1710 3540 1720 3700
rect 1780 3540 1790 3700
rect 2020 3540 2030 3700
rect 2090 3540 2100 3700
rect 2340 3540 2350 3700
rect 2410 3540 2420 3700
rect 2650 3540 2660 3700
rect 2720 3540 2730 3700
rect 280 3300 290 3460
rect 350 3300 360 3460
rect 600 3300 610 3460
rect 670 3300 680 3460
rect 920 3300 930 3460
rect 990 3300 1000 3460
rect 1230 3300 1240 3460
rect 1300 3300 1310 3460
rect 1550 3300 1560 3460
rect 1620 3300 1630 3460
rect 1860 3300 1870 3460
rect 1930 3300 1940 3460
rect 2180 3300 2190 3460
rect 2250 3300 2260 3460
rect 2500 3300 2510 3460
rect 2570 3300 2580 3460
rect 2760 3260 2860 3730
rect 0 3110 2860 3260
rect 0 2650 100 3110
rect 280 2920 290 3080
rect 350 2920 360 3080
rect 600 2920 610 3080
rect 670 2920 680 3080
rect 920 2920 930 3080
rect 990 2920 1000 3080
rect 1230 2920 1240 3080
rect 1300 2920 1310 3080
rect 1550 2920 1560 3080
rect 1620 2920 1630 3080
rect 1860 2920 1870 3080
rect 1930 2920 1940 3080
rect 2180 2920 2190 3080
rect 2250 2920 2260 3080
rect 2500 2920 2510 3080
rect 2570 2920 2580 3080
rect 130 2680 140 2840
rect 200 2680 210 2840
rect 440 2680 450 2840
rect 510 2680 520 2840
rect 760 2680 770 2840
rect 830 2680 840 2840
rect 1080 2680 1090 2840
rect 1150 2680 1160 2840
rect 1390 2680 1400 2840
rect 1460 2680 1470 2840
rect 1710 2680 1720 2840
rect 1780 2680 1790 2840
rect 2020 2680 2030 2840
rect 2090 2680 2100 2840
rect 2340 2680 2350 2840
rect 2410 2680 2420 2840
rect 2650 2680 2660 2840
rect 2720 2680 2730 2840
rect 2760 2650 2860 3110
rect 0 2500 2860 2650
rect 0 2030 100 2500
rect 130 2300 140 2460
rect 200 2300 210 2460
rect 440 2300 450 2460
rect 510 2300 520 2460
rect 760 2300 770 2460
rect 830 2300 840 2460
rect 1080 2300 1090 2460
rect 1150 2300 1160 2460
rect 1390 2300 1400 2460
rect 1460 2300 1470 2460
rect 1710 2300 1720 2460
rect 1780 2300 1790 2460
rect 2020 2300 2030 2460
rect 2090 2300 2100 2460
rect 2340 2300 2350 2460
rect 2410 2300 2420 2460
rect 2650 2300 2660 2460
rect 2720 2300 2730 2460
rect 280 2060 290 2220
rect 350 2060 360 2220
rect 600 2060 610 2220
rect 670 2060 680 2220
rect 920 2060 930 2220
rect 990 2060 1000 2220
rect 1230 2060 1240 2220
rect 1300 2060 1310 2220
rect 1550 2060 1560 2220
rect 1620 2060 1630 2220
rect 1860 2060 1870 2220
rect 1930 2060 1940 2220
rect 2180 2060 2190 2220
rect 2250 2060 2260 2220
rect 2500 2060 2510 2220
rect 2570 2060 2580 2220
rect 2760 2030 2860 2500
rect 0 1880 2860 2030
rect 0 1410 100 1880
rect 280 1690 290 1850
rect 350 1690 360 1850
rect 600 1690 610 1850
rect 670 1690 680 1850
rect 920 1690 930 1850
rect 990 1690 1000 1850
rect 1230 1690 1240 1850
rect 1300 1690 1310 1850
rect 1550 1690 1560 1850
rect 1620 1690 1630 1850
rect 1860 1690 1870 1850
rect 1930 1690 1940 1850
rect 2180 1690 2190 1850
rect 2250 1690 2260 1850
rect 2500 1690 2510 1850
rect 2570 1690 2580 1850
rect 130 1450 140 1610
rect 200 1450 210 1610
rect 440 1450 450 1610
rect 510 1450 520 1610
rect 760 1450 770 1610
rect 830 1450 840 1610
rect 1080 1450 1090 1610
rect 1150 1450 1160 1610
rect 1390 1450 1400 1610
rect 1460 1450 1470 1610
rect 1710 1450 1720 1610
rect 1780 1450 1790 1610
rect 2020 1450 2030 1610
rect 2090 1450 2100 1610
rect 2340 1450 2350 1610
rect 2410 1450 2420 1610
rect 2650 1450 2660 1610
rect 2720 1450 2730 1610
rect 2760 1410 2860 1880
rect 0 1260 2860 1410
rect 0 790 100 1260
rect 130 1070 140 1230
rect 200 1070 210 1230
rect 440 1070 450 1230
rect 510 1070 520 1230
rect 760 1070 770 1230
rect 830 1070 840 1230
rect 1080 1070 1090 1230
rect 1150 1070 1160 1230
rect 1390 1070 1400 1230
rect 1460 1070 1470 1230
rect 1710 1070 1720 1230
rect 1780 1070 1790 1230
rect 2020 1070 2030 1230
rect 2090 1070 2100 1230
rect 2340 1070 2350 1230
rect 2410 1070 2420 1230
rect 2650 1070 2660 1230
rect 2720 1070 2730 1230
rect 280 830 290 990
rect 350 830 360 990
rect 600 830 610 990
rect 670 830 680 990
rect 920 830 930 990
rect 990 830 1000 990
rect 1230 830 1240 990
rect 1300 830 1310 990
rect 1550 830 1560 990
rect 1620 830 1630 990
rect 1860 830 1870 990
rect 1930 830 1940 990
rect 2180 830 2190 990
rect 2250 830 2260 990
rect 2500 830 2510 990
rect 2570 830 2580 990
rect 2760 790 2860 1260
rect 0 640 2860 790
rect 0 180 100 640
rect 280 450 290 610
rect 350 450 360 610
rect 600 450 610 610
rect 670 450 680 610
rect 920 450 930 610
rect 990 450 1000 610
rect 1230 450 1240 610
rect 1300 450 1310 610
rect 1550 450 1560 610
rect 1620 450 1630 610
rect 1860 450 1870 610
rect 1930 450 1940 610
rect 2180 450 2190 610
rect 2250 450 2260 610
rect 2500 450 2510 610
rect 2570 450 2580 610
rect 130 210 140 370
rect 200 210 210 370
rect 440 210 450 370
rect 510 210 520 370
rect 760 210 770 370
rect 830 210 840 370
rect 1080 210 1090 370
rect 1150 210 1160 370
rect 1390 210 1400 370
rect 1460 210 1470 370
rect 1710 210 1720 370
rect 1780 210 1790 370
rect 2020 210 2030 370
rect 2090 210 2100 370
rect 2340 210 2350 370
rect 2410 210 2420 370
rect 2650 210 2660 370
rect 2720 210 2730 370
rect 2760 180 2860 640
rect 0 80 2860 180
rect 980 46 990 50
rect 978 -70 990 46
rect 1950 46 1960 50
rect 1950 -70 1962 46
rect 978 -76 1962 -70
<< via1 >>
rect 140 7460 200 7620
rect 330 7460 390 7620
rect 520 7460 580 7620
rect 710 7460 770 7620
rect 910 7460 970 7620
rect 1100 7460 1160 7620
rect 1290 7460 1350 7620
rect 1480 7460 1540 7620
rect 1670 7460 1730 7620
rect 230 7220 290 7380
rect 430 7220 490 7380
rect 620 7220 680 7380
rect 810 7220 870 7380
rect 1000 7220 1060 7380
rect 1190 7220 1250 7380
rect 1390 7220 1450 7380
rect 1580 7220 1640 7380
rect 230 6850 290 7010
rect 430 6850 490 7010
rect 620 6850 680 7010
rect 810 6850 870 7010
rect 1000 6850 1060 7010
rect 1190 6850 1250 7010
rect 1390 6850 1450 7010
rect 1580 6850 1640 7010
rect 140 6610 200 6770
rect 330 6610 390 6770
rect 520 6610 580 6770
rect 710 6610 770 6770
rect 910 6610 970 6770
rect 1100 6610 1160 6770
rect 1290 6610 1350 6770
rect 1480 6610 1540 6770
rect 1670 6610 1730 6770
rect 140 6230 200 6390
rect 330 6230 390 6390
rect 520 6230 580 6390
rect 710 6230 770 6390
rect 910 6230 970 6390
rect 1100 6230 1160 6390
rect 1290 6230 1350 6390
rect 1480 6230 1540 6390
rect 1670 6230 1730 6390
rect 230 5990 290 6150
rect 430 5990 490 6150
rect 620 5990 680 6150
rect 810 5990 870 6150
rect 1000 5990 1060 6150
rect 1190 5990 1250 6150
rect 1390 5990 1450 6150
rect 1580 5990 1640 6150
rect 230 5610 290 5770
rect 430 5610 490 5770
rect 620 5610 680 5770
rect 810 5610 870 5770
rect 1000 5610 1060 5770
rect 1190 5610 1250 5770
rect 1390 5610 1450 5770
rect 1580 5610 1640 5770
rect 140 5370 200 5530
rect 330 5370 390 5530
rect 520 5370 580 5530
rect 710 5370 770 5530
rect 910 5370 970 5530
rect 1100 5370 1160 5530
rect 1290 5370 1350 5530
rect 1480 5370 1540 5530
rect 1670 5370 1730 5530
rect 1020 5140 1730 5210
rect 140 4780 200 4940
rect 450 4780 510 4940
rect 770 4780 830 4940
rect 1090 4780 1150 4940
rect 1400 4780 1460 4940
rect 1720 4780 1780 4940
rect 2030 4780 2090 4940
rect 2350 4780 2410 4940
rect 2660 4780 2720 4940
rect 290 4540 350 4700
rect 610 4540 670 4700
rect 930 4540 990 4700
rect 1240 4540 1300 4700
rect 1560 4540 1620 4700
rect 1870 4540 1930 4700
rect 2190 4540 2250 4700
rect 2510 4540 2570 4700
rect 290 4160 350 4320
rect 610 4160 670 4320
rect 930 4160 990 4320
rect 1240 4160 1300 4320
rect 1560 4160 1620 4320
rect 1870 4160 1930 4320
rect 2190 4160 2250 4320
rect 2510 4160 2570 4320
rect 140 3920 200 4080
rect 450 3920 510 4080
rect 770 3920 830 4080
rect 1090 3920 1150 4080
rect 1400 3920 1460 4080
rect 1720 3920 1780 4080
rect 2030 3920 2090 4080
rect 2350 3920 2410 4080
rect 2660 3920 2720 4080
rect 140 3540 200 3700
rect 450 3540 510 3700
rect 770 3540 830 3700
rect 1090 3540 1150 3700
rect 1400 3540 1460 3700
rect 1720 3540 1780 3700
rect 2030 3540 2090 3700
rect 2350 3540 2410 3700
rect 2660 3540 2720 3700
rect 290 3300 350 3460
rect 610 3300 670 3460
rect 930 3300 990 3460
rect 1240 3300 1300 3460
rect 1560 3300 1620 3460
rect 1870 3300 1930 3460
rect 2190 3300 2250 3460
rect 2510 3300 2570 3460
rect 290 2920 350 3080
rect 610 2920 670 3080
rect 930 2920 990 3080
rect 1240 2920 1300 3080
rect 1560 2920 1620 3080
rect 1870 2920 1930 3080
rect 2190 2920 2250 3080
rect 2510 2920 2570 3080
rect 140 2680 200 2840
rect 450 2680 510 2840
rect 770 2680 830 2840
rect 1090 2680 1150 2840
rect 1400 2680 1460 2840
rect 1720 2680 1780 2840
rect 2030 2680 2090 2840
rect 2350 2680 2410 2840
rect 2660 2680 2720 2840
rect 140 2300 200 2460
rect 450 2300 510 2460
rect 770 2300 830 2460
rect 1090 2300 1150 2460
rect 1400 2300 1460 2460
rect 1720 2300 1780 2460
rect 2030 2300 2090 2460
rect 2350 2300 2410 2460
rect 2660 2300 2720 2460
rect 290 2060 350 2220
rect 610 2060 670 2220
rect 930 2060 990 2220
rect 1240 2060 1300 2220
rect 1560 2060 1620 2220
rect 1870 2060 1930 2220
rect 2190 2060 2250 2220
rect 2510 2060 2570 2220
rect 290 1690 350 1850
rect 610 1690 670 1850
rect 930 1690 990 1850
rect 1240 1690 1300 1850
rect 1560 1690 1620 1850
rect 1870 1690 1930 1850
rect 2190 1690 2250 1850
rect 2510 1690 2570 1850
rect 140 1450 200 1610
rect 450 1450 510 1610
rect 770 1450 830 1610
rect 1090 1450 1150 1610
rect 1400 1450 1460 1610
rect 1720 1450 1780 1610
rect 2030 1450 2090 1610
rect 2350 1450 2410 1610
rect 2660 1450 2720 1610
rect 140 1070 200 1230
rect 450 1070 510 1230
rect 770 1070 830 1230
rect 1090 1070 1150 1230
rect 1400 1070 1460 1230
rect 1720 1070 1780 1230
rect 2030 1070 2090 1230
rect 2350 1070 2410 1230
rect 2660 1070 2720 1230
rect 290 830 350 990
rect 610 830 670 990
rect 930 830 990 990
rect 1240 830 1300 990
rect 1560 830 1620 990
rect 1870 830 1930 990
rect 2190 830 2250 990
rect 2510 830 2570 990
rect 290 450 350 610
rect 610 450 670 610
rect 930 450 990 610
rect 1240 450 1300 610
rect 1560 450 1620 610
rect 1870 450 1930 610
rect 2190 450 2250 610
rect 2510 450 2570 610
rect 140 210 200 370
rect 450 210 510 370
rect 770 210 830 370
rect 1090 210 1150 370
rect 1400 210 1460 370
rect 1720 210 1780 370
rect 2030 210 2090 370
rect 2350 210 2410 370
rect 2660 210 2720 370
rect 990 40 1950 50
rect 990 -60 1950 40
<< metal2 >>
rect 140 7620 200 7630
rect 330 7620 390 7630
rect 520 7620 580 7630
rect 710 7620 770 7630
rect 910 7620 1730 7630
rect 200 7460 330 7620
rect 390 7460 520 7620
rect 580 7460 710 7620
rect 770 7460 910 7620
rect 970 7460 990 7620
rect 140 7450 200 7460
rect 330 7450 390 7460
rect 520 7450 580 7460
rect 710 7450 770 7460
rect 910 7450 1730 7460
rect 140 7380 870 7390
rect 1000 7380 1060 7390
rect 1190 7380 1250 7390
rect 1390 7380 1450 7390
rect 1580 7380 1640 7390
rect 870 7220 1000 7380
rect 1060 7220 1190 7380
rect 1250 7220 1390 7380
rect 1450 7220 1580 7380
rect 140 7210 870 7220
rect 1000 7210 1060 7220
rect 1190 7210 1250 7220
rect 1390 7210 1450 7220
rect 1580 7210 1640 7220
rect 140 7010 870 7020
rect 1000 7010 1060 7020
rect 1190 7010 1250 7020
rect 1390 7010 1450 7020
rect 1580 7010 1640 7020
rect 870 6850 1000 7010
rect 1060 6850 1190 7010
rect 1250 6850 1390 7010
rect 1450 6850 1580 7010
rect 140 6840 870 6850
rect 1000 6840 1060 6850
rect 1190 6840 1250 6850
rect 1390 6840 1450 6850
rect 1580 6840 1640 6850
rect 140 6770 200 6780
rect 330 6770 390 6780
rect 520 6770 580 6780
rect 710 6770 770 6780
rect 910 6770 1730 6780
rect 200 6610 330 6770
rect 390 6610 520 6770
rect 580 6610 710 6770
rect 770 6610 910 6770
rect 970 6610 990 6770
rect 140 6600 200 6610
rect 330 6600 390 6610
rect 520 6600 580 6610
rect 710 6600 770 6610
rect 910 6600 1730 6610
rect 140 6390 200 6400
rect 330 6390 390 6400
rect 520 6390 580 6400
rect 710 6390 770 6400
rect 910 6390 1730 6400
rect 200 6230 330 6390
rect 390 6230 520 6390
rect 580 6230 710 6390
rect 770 6230 910 6390
rect 970 6230 990 6390
rect 140 6220 200 6230
rect 330 6220 390 6230
rect 520 6220 580 6230
rect 710 6220 770 6230
rect 910 6220 1730 6230
rect 140 6150 870 6160
rect 1000 6150 1060 6160
rect 1190 6150 1250 6160
rect 1390 6150 1450 6160
rect 1580 6150 1640 6160
rect 870 5990 1000 6150
rect 1060 5990 1190 6150
rect 1250 5990 1390 6150
rect 1450 5990 1580 6150
rect 140 5980 870 5990
rect 1000 5980 1060 5990
rect 1190 5980 1250 5990
rect 1390 5980 1450 5990
rect 1580 5980 1640 5990
rect 140 5770 870 5780
rect 1000 5770 1060 5780
rect 1190 5770 1250 5780
rect 1390 5770 1450 5780
rect 1580 5770 1640 5780
rect 870 5610 1000 5770
rect 1060 5610 1190 5770
rect 1250 5610 1390 5770
rect 1450 5610 1580 5770
rect 140 5600 870 5610
rect 1000 5600 1060 5610
rect 1190 5600 1250 5610
rect 1390 5600 1450 5610
rect 1580 5600 1640 5610
rect 140 5530 200 5540
rect 330 5530 390 5540
rect 520 5530 580 5540
rect 710 5530 770 5540
rect 910 5530 1730 5540
rect 200 5370 330 5530
rect 390 5370 520 5530
rect 580 5370 710 5530
rect 770 5370 910 5530
rect 970 5370 990 5530
rect 140 5360 200 5370
rect 330 5360 390 5370
rect 520 5360 580 5370
rect 710 5360 770 5370
rect 910 5360 1730 5370
rect 1020 5210 1740 5230
rect 1730 5140 1740 5210
rect 1020 4950 1740 5140
rect 140 4940 200 4950
rect 450 4940 510 4950
rect 770 4940 830 4950
rect 1010 4940 1900 4950
rect 2030 4940 2090 4950
rect 2350 4940 2410 4950
rect 2660 4940 2720 4950
rect 200 4780 450 4940
rect 510 4780 770 4940
rect 830 4780 1010 4940
rect 1900 4780 2030 4940
rect 2090 4780 2350 4940
rect 2410 4780 2660 4940
rect 140 4770 200 4780
rect 450 4770 510 4780
rect 770 4770 830 4780
rect 1010 4770 1900 4780
rect 2030 4770 2090 4780
rect 2350 4770 2410 4780
rect 2660 4770 2720 4780
rect 140 4700 870 4710
rect 930 4700 990 4710
rect 1240 4700 1300 4710
rect 1560 4700 1620 4710
rect 1870 4700 1930 4710
rect 2190 4700 2250 4710
rect 2510 4700 2570 4710
rect 870 4540 930 4700
rect 990 4540 1240 4700
rect 1300 4540 1560 4700
rect 1620 4540 1870 4700
rect 1930 4540 2190 4700
rect 2250 4540 2510 4700
rect 140 4530 870 4540
rect 930 4530 990 4540
rect 1240 4530 1300 4540
rect 1560 4530 1620 4540
rect 1870 4530 1930 4540
rect 2190 4530 2250 4540
rect 2510 4530 2570 4540
rect 140 4320 870 4330
rect 930 4320 990 4330
rect 1240 4320 1300 4330
rect 1560 4320 1620 4330
rect 1870 4320 1930 4330
rect 2190 4320 2250 4330
rect 2510 4320 2570 4330
rect 870 4160 930 4320
rect 990 4160 1240 4320
rect 1300 4160 1560 4320
rect 1620 4160 1870 4320
rect 1930 4160 2190 4320
rect 2250 4160 2510 4320
rect 140 4150 870 4160
rect 930 4150 990 4160
rect 1240 4150 1300 4160
rect 1560 4150 1620 4160
rect 1870 4150 1930 4160
rect 2190 4150 2250 4160
rect 2510 4150 2570 4160
rect 140 4080 200 4090
rect 450 4080 510 4090
rect 770 4080 830 4090
rect 1010 4080 1900 4090
rect 2030 4080 2090 4090
rect 2350 4080 2410 4090
rect 2660 4080 2720 4090
rect 200 3920 450 4080
rect 510 3920 770 4080
rect 830 3920 1010 4080
rect 1900 3920 2030 4080
rect 2090 3920 2350 4080
rect 2410 3920 2660 4080
rect 140 3910 200 3920
rect 450 3910 510 3920
rect 770 3910 830 3920
rect 1010 3910 1900 3920
rect 2030 3910 2090 3920
rect 2350 3910 2410 3920
rect 2660 3910 2720 3920
rect 140 3700 200 3710
rect 450 3700 510 3710
rect 770 3700 830 3710
rect 1010 3700 1900 3710
rect 2030 3700 2090 3710
rect 2350 3700 2410 3710
rect 2660 3700 2720 3710
rect 200 3540 450 3700
rect 510 3540 770 3700
rect 830 3540 1010 3700
rect 1900 3540 2030 3700
rect 2090 3540 2350 3700
rect 2410 3540 2660 3700
rect 140 3530 200 3540
rect 450 3530 510 3540
rect 770 3530 830 3540
rect 1010 3530 1900 3540
rect 2030 3530 2090 3540
rect 2350 3530 2410 3540
rect 2660 3530 2720 3540
rect 140 3460 870 3470
rect 930 3460 990 3470
rect 1240 3460 1300 3470
rect 1560 3460 1620 3470
rect 1870 3460 1930 3470
rect 2190 3460 2250 3470
rect 2510 3460 2570 3470
rect 870 3300 930 3460
rect 990 3300 1240 3460
rect 1300 3300 1560 3460
rect 1620 3300 1870 3460
rect 1930 3300 2190 3460
rect 2250 3300 2510 3460
rect 140 3290 870 3300
rect 930 3290 990 3300
rect 1240 3290 1300 3300
rect 1560 3290 1620 3300
rect 1870 3290 1930 3300
rect 2190 3290 2250 3300
rect 2510 3290 2570 3300
rect 140 3080 870 3090
rect 930 3080 990 3090
rect 1240 3080 1300 3090
rect 1560 3080 1620 3090
rect 1870 3080 1930 3090
rect 2190 3080 2250 3090
rect 2510 3080 2570 3090
rect 870 2920 930 3080
rect 990 2920 1240 3080
rect 1300 2920 1560 3080
rect 1620 2920 1870 3080
rect 1930 2920 2190 3080
rect 2250 2920 2510 3080
rect 140 2910 870 2920
rect 930 2910 990 2920
rect 1240 2910 1300 2920
rect 1560 2910 1620 2920
rect 1870 2910 1930 2920
rect 2190 2910 2250 2920
rect 2510 2910 2570 2920
rect 140 2840 200 2850
rect 450 2840 510 2850
rect 770 2840 830 2850
rect 1010 2840 1900 2850
rect 2030 2840 2090 2850
rect 2350 2840 2410 2850
rect 2660 2840 2720 2850
rect 200 2680 450 2840
rect 510 2680 770 2840
rect 830 2680 1010 2840
rect 1900 2680 2030 2840
rect 2090 2680 2350 2840
rect 2410 2680 2660 2840
rect 140 2670 200 2680
rect 450 2670 510 2680
rect 770 2670 830 2680
rect 1010 2670 1900 2680
rect 2030 2670 2090 2680
rect 2350 2670 2410 2680
rect 2660 2670 2720 2680
rect 140 2460 200 2470
rect 450 2460 510 2470
rect 770 2460 830 2470
rect 1010 2460 1900 2470
rect 2030 2460 2090 2470
rect 2350 2460 2410 2470
rect 2660 2460 2720 2470
rect 200 2300 450 2460
rect 510 2300 770 2460
rect 830 2300 1010 2460
rect 1900 2300 2030 2460
rect 2090 2300 2350 2460
rect 2410 2300 2660 2460
rect 140 2290 200 2300
rect 450 2290 510 2300
rect 770 2290 830 2300
rect 1010 2290 1900 2300
rect 2030 2290 2090 2300
rect 2350 2290 2410 2300
rect 2660 2290 2720 2300
rect 140 2220 870 2230
rect 930 2220 990 2230
rect 1240 2220 1300 2230
rect 1560 2220 1620 2230
rect 1870 2220 1930 2230
rect 2190 2220 2250 2230
rect 2510 2220 2570 2230
rect 870 2060 930 2220
rect 990 2060 1240 2220
rect 1300 2060 1560 2220
rect 1620 2060 1870 2220
rect 1930 2060 2190 2220
rect 2250 2060 2510 2220
rect 140 2050 870 2060
rect 930 2050 990 2060
rect 1240 2050 1300 2060
rect 1560 2050 1620 2060
rect 1870 2050 1930 2060
rect 2190 2050 2250 2060
rect 2510 2050 2570 2060
rect 140 1850 870 1860
rect 930 1850 990 1860
rect 1240 1850 1300 1860
rect 1560 1850 1620 1860
rect 1870 1850 1930 1860
rect 2190 1850 2250 1860
rect 2510 1850 2570 1860
rect 870 1690 930 1850
rect 990 1690 1240 1850
rect 1300 1690 1560 1850
rect 1620 1690 1870 1850
rect 1930 1690 2190 1850
rect 2250 1690 2510 1850
rect 140 1680 870 1690
rect 930 1680 990 1690
rect 1240 1680 1300 1690
rect 1560 1680 1620 1690
rect 1870 1680 1930 1690
rect 2190 1680 2250 1690
rect 2510 1680 2570 1690
rect 140 1610 200 1620
rect 450 1610 510 1620
rect 770 1610 830 1620
rect 1010 1610 1900 1620
rect 2030 1610 2090 1620
rect 2350 1610 2410 1620
rect 2660 1610 2720 1620
rect 200 1450 450 1610
rect 510 1450 770 1610
rect 830 1450 1010 1610
rect 1900 1450 2030 1610
rect 2090 1450 2350 1610
rect 2410 1450 2660 1610
rect 140 1440 200 1450
rect 450 1440 510 1450
rect 770 1440 830 1450
rect 1010 1440 1900 1450
rect 2030 1440 2090 1450
rect 2350 1440 2410 1450
rect 2660 1440 2720 1450
rect 140 1230 200 1240
rect 450 1230 510 1240
rect 770 1230 830 1240
rect 1010 1230 1900 1240
rect 2030 1230 2090 1240
rect 2350 1230 2410 1240
rect 2660 1230 2720 1240
rect 200 1070 450 1230
rect 510 1070 770 1230
rect 830 1070 1010 1230
rect 1900 1070 2030 1230
rect 2090 1070 2350 1230
rect 2410 1070 2660 1230
rect 140 1060 200 1070
rect 450 1060 510 1070
rect 770 1060 830 1070
rect 1010 1060 1900 1070
rect 2030 1060 2090 1070
rect 2350 1060 2410 1070
rect 2660 1060 2720 1070
rect 140 990 870 1000
rect 930 990 990 1000
rect 1240 990 1300 1000
rect 1560 990 1620 1000
rect 1870 990 1930 1000
rect 2190 990 2250 1000
rect 2510 990 2570 1000
rect 870 830 930 990
rect 990 830 1240 990
rect 1300 830 1560 990
rect 1620 830 1870 990
rect 1930 830 2190 990
rect 2250 830 2510 990
rect 140 820 870 830
rect 930 820 990 830
rect 1240 820 1300 830
rect 1560 820 1620 830
rect 1870 820 1930 830
rect 2190 820 2250 830
rect 2510 820 2570 830
rect 140 610 870 620
rect 930 610 990 620
rect 1240 610 1300 620
rect 1560 610 1620 620
rect 1870 610 1930 620
rect 2190 610 2250 620
rect 2510 610 2570 620
rect 870 450 930 610
rect 990 450 1240 610
rect 1300 450 1560 610
rect 1620 450 1870 610
rect 1930 450 2190 610
rect 2250 450 2510 610
rect 140 440 870 450
rect 930 440 990 450
rect 1240 440 1300 450
rect 1560 440 1620 450
rect 1870 440 1930 450
rect 2190 440 2250 450
rect 2510 440 2570 450
rect 140 370 200 380
rect 450 370 510 380
rect 770 370 830 380
rect 1010 370 1900 380
rect 2030 370 2090 380
rect 2350 370 2410 380
rect 2660 370 2720 380
rect 200 210 450 370
rect 510 210 770 370
rect 830 210 1010 370
rect 1900 210 2030 370
rect 2090 210 2350 370
rect 2410 210 2660 370
rect 140 200 200 210
rect 450 200 510 210
rect 770 200 830 210
rect 990 50 1950 210
rect 2030 200 2090 210
rect 2350 200 2410 210
rect 2660 200 2720 210
rect 990 -70 1950 -60
<< via2 >>
rect 990 7460 1100 7620
rect 1100 7460 1160 7620
rect 1160 7460 1290 7620
rect 1290 7460 1350 7620
rect 1350 7460 1480 7620
rect 1480 7460 1540 7620
rect 1540 7460 1670 7620
rect 1670 7460 1730 7620
rect 140 7220 230 7380
rect 230 7220 290 7380
rect 290 7220 430 7380
rect 430 7220 490 7380
rect 490 7220 620 7380
rect 620 7220 680 7380
rect 680 7220 810 7380
rect 810 7220 870 7380
rect 140 6850 230 7010
rect 230 6850 290 7010
rect 290 6850 430 7010
rect 430 6850 490 7010
rect 490 6850 620 7010
rect 620 6850 680 7010
rect 680 6850 810 7010
rect 810 6850 870 7010
rect 990 6610 1100 6770
rect 1100 6610 1160 6770
rect 1160 6610 1290 6770
rect 1290 6610 1350 6770
rect 1350 6610 1480 6770
rect 1480 6610 1540 6770
rect 1540 6610 1670 6770
rect 1670 6610 1730 6770
rect 990 6230 1100 6390
rect 1100 6230 1160 6390
rect 1160 6230 1290 6390
rect 1290 6230 1350 6390
rect 1350 6230 1480 6390
rect 1480 6230 1540 6390
rect 1540 6230 1670 6390
rect 1670 6230 1730 6390
rect 140 5990 230 6150
rect 230 5990 290 6150
rect 290 5990 430 6150
rect 430 5990 490 6150
rect 490 5990 620 6150
rect 620 5990 680 6150
rect 680 5990 810 6150
rect 810 5990 870 6150
rect 140 5610 230 5770
rect 230 5610 290 5770
rect 290 5610 430 5770
rect 430 5610 490 5770
rect 490 5610 620 5770
rect 620 5610 680 5770
rect 680 5610 810 5770
rect 810 5610 870 5770
rect 990 5370 1100 5530
rect 1100 5370 1160 5530
rect 1160 5370 1290 5530
rect 1290 5370 1350 5530
rect 1350 5370 1480 5530
rect 1480 5370 1540 5530
rect 1540 5370 1670 5530
rect 1670 5370 1730 5530
rect 1010 4780 1090 4940
rect 1090 4780 1150 4940
rect 1150 4780 1400 4940
rect 1400 4780 1460 4940
rect 1460 4780 1720 4940
rect 1720 4780 1780 4940
rect 1780 4780 1900 4940
rect 140 4540 290 4700
rect 290 4540 350 4700
rect 350 4540 610 4700
rect 610 4540 670 4700
rect 670 4540 870 4700
rect 140 4160 290 4320
rect 290 4160 350 4320
rect 350 4160 610 4320
rect 610 4160 670 4320
rect 670 4160 870 4320
rect 1010 3920 1090 4080
rect 1090 3920 1150 4080
rect 1150 3920 1400 4080
rect 1400 3920 1460 4080
rect 1460 3920 1720 4080
rect 1720 3920 1780 4080
rect 1780 3920 1900 4080
rect 1010 3540 1090 3700
rect 1090 3540 1150 3700
rect 1150 3540 1400 3700
rect 1400 3540 1460 3700
rect 1460 3540 1720 3700
rect 1720 3540 1780 3700
rect 1780 3540 1900 3700
rect 140 3300 290 3460
rect 290 3300 350 3460
rect 350 3300 610 3460
rect 610 3300 670 3460
rect 670 3300 870 3460
rect 140 2920 290 3080
rect 290 2920 350 3080
rect 350 2920 610 3080
rect 610 2920 670 3080
rect 670 2920 870 3080
rect 1010 2680 1090 2840
rect 1090 2680 1150 2840
rect 1150 2680 1400 2840
rect 1400 2680 1460 2840
rect 1460 2680 1720 2840
rect 1720 2680 1780 2840
rect 1780 2680 1900 2840
rect 1010 2300 1090 2460
rect 1090 2300 1150 2460
rect 1150 2300 1400 2460
rect 1400 2300 1460 2460
rect 1460 2300 1720 2460
rect 1720 2300 1780 2460
rect 1780 2300 1900 2460
rect 140 2060 290 2220
rect 290 2060 350 2220
rect 350 2060 610 2220
rect 610 2060 670 2220
rect 670 2060 870 2220
rect 140 1690 290 1850
rect 290 1690 350 1850
rect 350 1690 610 1850
rect 610 1690 670 1850
rect 670 1690 870 1850
rect 1010 1450 1090 1610
rect 1090 1450 1150 1610
rect 1150 1450 1400 1610
rect 1400 1450 1460 1610
rect 1460 1450 1720 1610
rect 1720 1450 1780 1610
rect 1780 1450 1900 1610
rect 1010 1070 1090 1230
rect 1090 1070 1150 1230
rect 1150 1070 1400 1230
rect 1400 1070 1460 1230
rect 1460 1070 1720 1230
rect 1720 1070 1780 1230
rect 1780 1070 1900 1230
rect 140 830 290 990
rect 290 830 350 990
rect 350 830 610 990
rect 610 830 670 990
rect 670 830 870 990
rect 140 450 290 610
rect 290 450 350 610
rect 350 450 610 610
rect 610 450 670 610
rect 670 450 870 610
rect 1010 210 1090 370
rect 1090 210 1150 370
rect 1150 210 1400 370
rect 1400 210 1460 370
rect 1460 210 1720 370
rect 1720 210 1780 370
rect 1780 210 1900 370
<< metal3 >>
rect 990 7625 1730 7840
rect 980 7620 1740 7625
rect 980 7460 990 7620
rect 1730 7460 1740 7620
rect 980 7455 1740 7460
rect 140 7385 870 7390
rect 130 7380 880 7385
rect 130 7220 140 7380
rect 870 7220 880 7380
rect 130 7215 880 7220
rect 140 7015 870 7215
rect 130 7010 880 7015
rect 130 6850 140 7010
rect 870 6850 880 7010
rect 130 6845 880 6850
rect 140 6155 870 6845
rect 990 6775 1730 7455
rect 980 6770 1740 6775
rect 980 6610 990 6770
rect 1730 6610 1740 6770
rect 980 6605 1740 6610
rect 990 6395 1730 6605
rect 980 6390 1740 6395
rect 980 6230 990 6390
rect 1730 6230 1740 6390
rect 980 6225 1740 6230
rect 130 6150 880 6155
rect 130 5990 140 6150
rect 870 5990 880 6150
rect 130 5985 880 5990
rect 140 5775 870 5985
rect 130 5770 880 5775
rect 130 5610 140 5770
rect 870 5610 880 5770
rect 130 5605 880 5610
rect 140 4705 870 5605
rect 990 5535 1730 6225
rect 980 5530 1740 5535
rect 980 5370 990 5530
rect 1730 5370 1740 5530
rect 980 5365 1740 5370
rect 1000 4940 1910 4945
rect 1000 4780 1010 4940
rect 1900 4780 1910 4940
rect 1000 4775 1910 4780
rect 130 4700 880 4705
rect 130 4540 140 4700
rect 870 4540 880 4700
rect 130 4535 880 4540
rect 140 4325 870 4535
rect 130 4320 880 4325
rect 130 4160 140 4320
rect 870 4160 880 4320
rect 130 4155 880 4160
rect 140 3465 870 4155
rect 1010 4085 1900 4775
rect 1000 4080 1910 4085
rect 1000 3920 1010 4080
rect 1900 3920 1910 4080
rect 1000 3915 1910 3920
rect 1010 3705 1900 3915
rect 1000 3700 1910 3705
rect 1000 3540 1010 3700
rect 1900 3540 1910 3700
rect 1000 3535 1910 3540
rect 130 3460 880 3465
rect 130 3300 140 3460
rect 870 3300 880 3460
rect 130 3295 880 3300
rect 140 3085 870 3295
rect 130 3080 880 3085
rect 130 2920 140 3080
rect 870 2920 880 3080
rect 130 2915 880 2920
rect 140 2225 870 2915
rect 1010 2845 1900 3535
rect 1000 2840 1910 2845
rect 1000 2680 1010 2840
rect 1900 2680 1910 2840
rect 1000 2675 1910 2680
rect 1010 2465 1900 2675
rect 1000 2460 1910 2465
rect 1000 2300 1010 2460
rect 1900 2300 1910 2460
rect 1000 2295 1910 2300
rect 130 2220 880 2225
rect 130 2060 140 2220
rect 870 2060 880 2220
rect 130 2055 880 2060
rect 140 1855 870 2055
rect 130 1850 880 1855
rect 130 1690 140 1850
rect 870 1690 880 1850
rect 130 1685 880 1690
rect 140 995 870 1685
rect 1010 1615 1900 2295
rect 1000 1610 1910 1615
rect 1000 1450 1010 1610
rect 1900 1450 1910 1610
rect 1000 1445 1910 1450
rect 1010 1235 1900 1445
rect 1000 1230 1910 1235
rect 1000 1070 1010 1230
rect 1900 1070 1910 1230
rect 1000 1065 1910 1070
rect 130 990 880 995
rect 130 830 140 990
rect 870 830 880 990
rect 130 825 880 830
rect 140 615 870 825
rect 130 610 880 615
rect 130 450 140 610
rect 870 450 880 610
rect 130 445 880 450
rect 1010 375 1900 1065
rect 1000 370 1910 375
rect 1000 210 1010 370
rect 1900 210 1910 370
rect 1000 205 1910 210
use outd_cmirror_transistors  outd_cmirror_transistors_0
timestamp 1647254192
transform 1 0 180 0 1 5340
box -180 -5340 2682 2494
<< end >>
