magic
tech sky130A
magscale 1 2
timestamp 1646042961
<< nwell >>
rect -2173 -618 -1507 618
rect -1253 -618 -587 618
rect -333 -618 333 618
rect 587 -618 1253 618
rect 1507 -618 2173 618
<< pwell >>
rect -2283 618 2283 728
rect -2283 -618 -2173 618
rect -1507 -618 -1253 618
rect -587 -618 -333 618
rect 333 -618 587 618
rect 1253 -618 1507 618
rect 2173 -618 2283 618
rect -2283 -728 2283 -618
<< varactor >>
rect -2040 -500 -1640 500
rect -1120 -500 -720 500
rect -200 -500 200 500
rect 720 -500 1120 500
rect 1640 -500 2040 500
<< psubdiff >>
rect -2247 658 -2151 692
rect 2151 658 2247 692
rect -2247 569 -2213 658
rect 2213 569 2247 658
rect -2247 -658 -2213 -569
rect 2213 -658 2247 -569
rect -2247 -692 -2124 -658
rect 2124 -692 2247 -658
<< nsubdiff >>
rect -2137 476 -2040 500
rect -2137 -476 -2125 476
rect -2091 -476 -2040 476
rect -2137 -500 -2040 -476
rect -1640 476 -1543 500
rect -1640 -476 -1589 476
rect -1555 -476 -1543 476
rect -1640 -500 -1543 -476
rect -1217 476 -1120 500
rect -1217 -476 -1205 476
rect -1171 -476 -1120 476
rect -1217 -500 -1120 -476
rect -720 476 -623 500
rect -720 -476 -669 476
rect -635 -476 -623 476
rect -720 -500 -623 -476
rect -297 476 -200 500
rect -297 -476 -285 476
rect -251 -476 -200 476
rect -297 -500 -200 -476
rect 200 476 297 500
rect 200 -476 251 476
rect 285 -476 297 476
rect 200 -500 297 -476
rect 623 476 720 500
rect 623 -476 635 476
rect 669 -476 720 476
rect 623 -500 720 -476
rect 1120 476 1217 500
rect 1120 -476 1171 476
rect 1205 -476 1217 476
rect 1120 -500 1217 -476
rect 1543 476 1640 500
rect 1543 -476 1555 476
rect 1589 -476 1640 476
rect 1543 -500 1640 -476
rect 2040 476 2137 500
rect 2040 -476 2091 476
rect 2125 -476 2137 476
rect 2040 -500 2137 -476
<< psubdiffcont >>
rect -2151 658 2151 692
rect -2247 -569 -2213 569
rect 2213 -569 2247 569
rect -2124 -692 2124 -658
<< nsubdiffcont >>
rect -2125 -476 -2091 476
rect -1589 -476 -1555 476
rect -1205 -476 -1171 476
rect -669 -476 -635 476
rect -285 -476 -251 476
rect 251 -476 285 476
rect 635 -476 669 476
rect 1171 -476 1205 476
rect 1555 -476 1589 476
rect 2091 -476 2125 476
<< poly >>
rect -2040 572 -1640 588
rect -2040 538 -2024 572
rect -1656 538 -1640 572
rect -2040 500 -1640 538
rect -1120 572 -720 588
rect -1120 538 -1104 572
rect -736 538 -720 572
rect -1120 500 -720 538
rect -200 572 200 588
rect -200 538 -184 572
rect 184 538 200 572
rect -200 500 200 538
rect 720 572 1120 588
rect 720 538 736 572
rect 1104 538 1120 572
rect 720 500 1120 538
rect 1640 572 2040 588
rect 1640 538 1656 572
rect 2024 538 2040 572
rect 1640 500 2040 538
rect -2040 -538 -1640 -500
rect -2040 -572 -2024 -538
rect -1656 -572 -1640 -538
rect -2040 -588 -1640 -572
rect -1120 -538 -720 -500
rect -1120 -572 -1104 -538
rect -736 -572 -720 -538
rect -1120 -588 -720 -572
rect -200 -538 200 -500
rect -200 -572 -184 -538
rect 184 -572 200 -538
rect -200 -588 200 -572
rect 720 -538 1120 -500
rect 720 -572 736 -538
rect 1104 -572 1120 -538
rect 720 -588 1120 -572
rect 1640 -538 2040 -500
rect 1640 -572 1656 -538
rect 2024 -572 2040 -538
rect 1640 -588 2040 -572
<< polycont >>
rect -2024 538 -1656 572
rect -1104 538 -736 572
rect -184 538 184 572
rect 736 538 1104 572
rect 1656 538 2024 572
rect -2024 -572 -1656 -538
rect -1104 -572 -736 -538
rect -184 -572 184 -538
rect 736 -572 1104 -538
rect 1656 -572 2024 -538
<< locali >>
rect -2247 658 -2151 692
rect 2151 658 2247 692
rect -2247 569 -2213 658
rect -2040 538 -2024 572
rect -1656 538 -1640 572
rect -1120 538 -1104 572
rect -736 538 -720 572
rect -200 538 -184 572
rect 184 538 200 572
rect 720 538 736 572
rect 1104 538 1120 572
rect 1640 538 1656 572
rect 2024 538 2040 572
rect 2213 569 2247 658
rect -2125 476 -2091 492
rect -2125 -492 -2091 -476
rect -1589 476 -1555 492
rect -1589 -492 -1555 -476
rect -1205 476 -1171 492
rect -1205 -492 -1171 -476
rect -669 476 -635 492
rect -669 -492 -635 -476
rect -285 476 -251 492
rect -285 -492 -251 -476
rect 251 476 285 492
rect 251 -492 285 -476
rect 635 476 669 492
rect 635 -492 669 -476
rect 1171 476 1205 492
rect 1171 -492 1205 -476
rect 1555 476 1589 492
rect 1555 -492 1589 -476
rect 2091 476 2125 492
rect 2091 -492 2125 -476
rect -2247 -658 -2213 -569
rect -2040 -572 -2024 -538
rect -1656 -572 -1640 -538
rect -1120 -572 -1104 -538
rect -736 -572 -720 -538
rect -200 -572 -184 -538
rect 184 -572 200 -538
rect 720 -572 736 -538
rect 1104 -572 1120 -538
rect 1640 -572 1656 -538
rect 2024 -572 2040 -538
rect 2213 -658 2247 -569
rect -2247 -692 -2124 -658
rect 2124 -692 2247 -658
<< viali >>
rect -2024 538 -1656 572
rect -1104 538 -736 572
rect -184 538 184 572
rect 736 538 1104 572
rect 1656 538 2024 572
rect -2125 -476 -2091 476
rect -1589 -476 -1555 476
rect -1205 -476 -1171 476
rect -669 -476 -635 476
rect -285 -476 -251 476
rect 251 -476 285 476
rect 635 -476 669 476
rect 1171 -476 1205 476
rect 1555 -476 1589 476
rect 2091 -476 2125 476
rect -2024 -572 -1656 -538
rect -1104 -572 -736 -538
rect -184 -572 184 -538
rect 736 -572 1104 -538
rect 1656 -572 2024 -538
<< metal1 >>
rect -2036 572 -1644 578
rect -2036 538 -2024 572
rect -1656 538 -1644 572
rect -2036 532 -1644 538
rect -1116 572 -724 578
rect -1116 538 -1104 572
rect -736 538 -724 572
rect -1116 532 -724 538
rect -196 572 196 578
rect -196 538 -184 572
rect 184 538 196 572
rect -196 532 196 538
rect 724 572 1116 578
rect 724 538 736 572
rect 1104 538 1116 572
rect 724 532 1116 538
rect 1644 572 2036 578
rect 1644 538 1656 572
rect 2024 538 2036 572
rect 1644 532 2036 538
rect -2131 476 -2085 488
rect -2131 -476 -2125 476
rect -2091 -476 -2085 476
rect -2131 -488 -2085 -476
rect -1595 476 -1549 488
rect -1595 -476 -1589 476
rect -1555 -476 -1549 476
rect -1595 -488 -1549 -476
rect -1211 476 -1165 488
rect -1211 -476 -1205 476
rect -1171 -476 -1165 476
rect -1211 -488 -1165 -476
rect -675 476 -629 488
rect -675 -476 -669 476
rect -635 -476 -629 476
rect -675 -488 -629 -476
rect -291 476 -245 488
rect -291 -476 -285 476
rect -251 -476 -245 476
rect -291 -488 -245 -476
rect 245 476 291 488
rect 245 -476 251 476
rect 285 -476 291 476
rect 245 -488 291 -476
rect 629 476 675 488
rect 629 -476 635 476
rect 669 -476 675 476
rect 629 -488 675 -476
rect 1165 476 1211 488
rect 1165 -476 1171 476
rect 1205 -476 1211 476
rect 1165 -488 1211 -476
rect 1549 476 1595 488
rect 1549 -476 1555 476
rect 1589 -476 1595 476
rect 1549 -488 1595 -476
rect 2085 476 2131 488
rect 2085 -476 2091 476
rect 2125 -476 2131 476
rect 2085 -488 2131 -476
rect -2036 -538 -1644 -532
rect -2036 -572 -2024 -538
rect -1656 -572 -1644 -538
rect -2036 -578 -1644 -572
rect -1116 -538 -724 -532
rect -1116 -572 -1104 -538
rect -736 -572 -724 -538
rect -1116 -578 -724 -572
rect -196 -538 196 -532
rect -196 -572 -184 -538
rect 184 -572 196 -538
rect -196 -578 196 -572
rect 724 -538 1116 -532
rect 724 -572 736 -538
rect 1104 -572 1116 -538
rect 724 -578 1116 -572
rect 1644 -538 2036 -532
rect 1644 -572 1656 -538
rect 2024 -572 2036 -538
rect 1644 -578 2036 -572
<< properties >>
string FIXED_BBOX -2230 -648 2230 648
string gencell sky130_fd_pr__cap_var_lvt
string library sky130
string parameters w 5 l 2 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.18 wmin 1.0 compatible {sky130_fd_pr__cap_var_lvt  sky130_fd_pr__cap_var_hvt sky130_fd_pr__cap_var} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
