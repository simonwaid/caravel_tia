magic
tech sky130A
magscale 1 2
timestamp 1647254192
<< pwell >>
rect -2683 -610 2683 610
<< nmos >>
rect -2487 -400 -1287 400
rect -1229 -400 -29 400
rect 29 -400 1229 400
rect 1287 -400 2487 400
<< ndiff >>
rect -2545 388 -2487 400
rect -2545 -388 -2533 388
rect -2499 -388 -2487 388
rect -2545 -400 -2487 -388
rect -1287 388 -1229 400
rect -1287 -388 -1275 388
rect -1241 -388 -1229 388
rect -1287 -400 -1229 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 1229 388 1287 400
rect 1229 -388 1241 388
rect 1275 -388 1287 388
rect 1229 -400 1287 -388
rect 2487 388 2545 400
rect 2487 -388 2499 388
rect 2533 -388 2545 388
rect 2487 -400 2545 -388
<< ndiffc >>
rect -2533 -388 -2499 388
rect -1275 -388 -1241 388
rect -17 -388 17 388
rect 1241 -388 1275 388
rect 2499 -388 2533 388
<< psubdiff >>
rect -2647 540 -2551 574
rect 2551 540 2647 574
rect -2647 478 -2613 540
rect 2613 478 2647 540
rect -2647 -540 -2613 -478
rect 2613 -540 2647 -478
rect -2647 -574 -2551 -540
rect 2551 -574 2647 -540
<< psubdiffcont >>
rect -2551 540 2551 574
rect -2647 -478 -2613 478
rect 2613 -478 2647 478
rect -2551 -574 2551 -540
<< poly >>
rect -2487 472 -1287 488
rect -2487 438 -2471 472
rect -1303 438 -1287 472
rect -2487 400 -1287 438
rect -1229 472 -29 488
rect -1229 438 -1213 472
rect -45 438 -29 472
rect -1229 400 -29 438
rect 29 472 1229 488
rect 29 438 45 472
rect 1213 438 1229 472
rect 29 400 1229 438
rect 1287 472 2487 488
rect 1287 438 1303 472
rect 2471 438 2487 472
rect 1287 400 2487 438
rect -2487 -438 -1287 -400
rect -2487 -472 -2471 -438
rect -1303 -472 -1287 -438
rect -2487 -488 -1287 -472
rect -1229 -438 -29 -400
rect -1229 -472 -1213 -438
rect -45 -472 -29 -438
rect -1229 -488 -29 -472
rect 29 -438 1229 -400
rect 29 -472 45 -438
rect 1213 -472 1229 -438
rect 29 -488 1229 -472
rect 1287 -438 2487 -400
rect 1287 -472 1303 -438
rect 2471 -472 2487 -438
rect 1287 -488 2487 -472
<< polycont >>
rect -2471 438 -1303 472
rect -1213 438 -45 472
rect 45 438 1213 472
rect 1303 438 2471 472
rect -2471 -472 -1303 -438
rect -1213 -472 -45 -438
rect 45 -472 1213 -438
rect 1303 -472 2471 -438
<< locali >>
rect -2647 540 -2551 574
rect 2551 540 2647 574
rect -2647 478 -2613 540
rect 2613 478 2647 540
rect -2487 438 -2471 472
rect -1303 438 -1287 472
rect -1229 438 -1213 472
rect -45 438 -29 472
rect 29 438 45 472
rect 1213 438 1229 472
rect 1287 438 1303 472
rect 2471 438 2487 472
rect -2533 388 -2499 404
rect -2533 -404 -2499 -388
rect -1275 388 -1241 404
rect -1275 -404 -1241 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 1241 388 1275 404
rect 1241 -404 1275 -388
rect 2499 388 2533 404
rect 2499 -404 2533 -388
rect -2487 -472 -2471 -438
rect -1303 -472 -1287 -438
rect -1229 -472 -1213 -438
rect -45 -472 -29 -438
rect 29 -472 45 -438
rect 1213 -472 1229 -438
rect 1287 -472 1303 -438
rect 2471 -472 2487 -438
rect -2647 -540 -2613 -478
rect 2613 -540 2647 -478
rect -2647 -574 -2551 -540
rect 2551 -574 2647 -540
<< viali >>
rect -2471 438 -1303 472
rect -1213 438 -45 472
rect 45 438 1213 472
rect 1303 438 2471 472
rect -2533 -388 -2499 388
rect -1275 -388 -1241 388
rect -17 -388 17 388
rect 1241 -388 1275 388
rect 2499 -388 2533 388
rect -2471 -472 -1303 -438
rect -1213 -472 -45 -438
rect 45 -472 1213 -438
rect 1303 -472 2471 -438
<< metal1 >>
rect -2483 472 -1291 478
rect -2483 438 -2471 472
rect -1303 438 -1291 472
rect -2483 432 -1291 438
rect -1225 472 -33 478
rect -1225 438 -1213 472
rect -45 438 -33 472
rect -1225 432 -33 438
rect 33 472 1225 478
rect 33 438 45 472
rect 1213 438 1225 472
rect 33 432 1225 438
rect 1291 472 2483 478
rect 1291 438 1303 472
rect 2471 438 2483 472
rect 1291 432 2483 438
rect -2539 388 -2493 400
rect -2539 -388 -2533 388
rect -2499 -388 -2493 388
rect -2539 -400 -2493 -388
rect -1281 388 -1235 400
rect -1281 -388 -1275 388
rect -1241 -388 -1235 388
rect -1281 -400 -1235 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 1235 388 1281 400
rect 1235 -388 1241 388
rect 1275 -388 1281 388
rect 1235 -400 1281 -388
rect 2493 388 2539 400
rect 2493 -388 2499 388
rect 2533 -388 2539 388
rect 2493 -400 2539 -388
rect -2483 -438 -1291 -432
rect -2483 -472 -2471 -438
rect -1303 -472 -1291 -438
rect -2483 -478 -1291 -472
rect -1225 -438 -33 -432
rect -1225 -472 -1213 -438
rect -45 -472 -33 -438
rect -1225 -478 -33 -472
rect 33 -438 1225 -432
rect 33 -472 45 -438
rect 1213 -472 1225 -438
rect 33 -478 1225 -472
rect 1291 -438 2483 -432
rect 1291 -472 1303 -438
rect 2471 -472 2483 -438
rect 1291 -478 2483 -472
<< properties >>
string FIXED_BBOX -2630 -557 2630 557
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 4 l 6 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
