magic
tech sky130A
magscale 1 2
timestamp 1645630008
<< locali >>
rect 17180 12710 22720 13000
rect 4360 12650 22720 12710
rect 4360 12600 22840 12650
rect 23190 12600 23240 13000
rect 4360 12590 17410 12600
rect 17170 11940 17410 12590
rect 17170 11700 17300 11940
rect 17400 11700 17410 11940
rect 17170 11470 17410 11700
rect 22680 11480 22840 12600
<< viali >>
rect 17300 11700 17400 11940
<< metal1 >>
rect 16760 13700 17860 13860
rect 16760 12820 16980 13700
rect 17680 13200 17860 13700
rect 17680 13000 17700 13200
rect 17840 13000 17860 13200
rect 17680 12980 17860 13000
rect 20980 12880 21160 15060
rect 22820 13360 23120 13380
rect 22820 13180 22840 13360
rect 23100 13180 23120 13360
rect 16760 12480 17020 12820
rect 20970 12680 20980 12880
rect 21160 12680 21170 12880
rect 16760 11560 16980 12480
rect 17294 11940 17406 11952
rect 17290 11700 17300 11940
rect 17400 11700 17410 11940
rect 17470 11700 17480 11940
rect 17560 11700 17570 11940
rect 17294 11688 17406 11700
rect 17600 11580 17800 12520
rect 18740 12488 18830 12522
rect 19998 12488 20088 12522
rect 21256 12488 21346 12522
rect 18730 12160 18740 12400
rect 18820 12160 18830 12400
rect 21250 12160 21260 12400
rect 21340 12160 21350 12400
rect 19990 11700 20000 11940
rect 20080 11700 20090 11940
rect 22510 11700 22520 11940
rect 22600 11700 22610 11940
rect 18740 11578 18830 11612
rect 19998 11578 20088 11612
rect 21256 11578 21346 11612
rect 22820 11580 23120 13180
rect 23460 11560 24300 12020
rect 24520 11560 25360 12020
rect 22920 9140 23760 9600
rect 24000 9140 24840 9600
rect 25050 9160 25060 9580
rect 25360 9160 25370 9580
<< via1 >>
rect 17700 13000 17840 13200
rect 22840 13180 23100 13360
rect 20980 12680 21160 12880
rect 17300 11700 17400 11940
rect 17480 11700 17560 11940
rect 18740 12160 18820 12400
rect 21260 12160 21340 12400
rect 20000 11700 20080 11940
rect 22520 11700 22600 11940
rect 25060 9160 25360 9580
<< metal2 >>
rect 16960 13630 17520 13680
rect 16680 13620 17520 13630
rect 17000 13480 17520 13620
rect 16680 13470 17520 13480
rect 16960 13420 17520 13470
rect 16680 12400 17100 13080
rect 17260 12880 17520 13420
rect 20900 13360 21120 13840
rect 17700 13200 17840 13210
rect 20900 13200 20920 13360
rect 17840 13100 20920 13200
rect 22840 13360 23100 13370
rect 22840 13170 23100 13180
rect 17840 13000 21120 13100
rect 17700 12990 17840 13000
rect 20980 12880 21160 12890
rect 23140 12880 23360 13700
rect 17260 12680 20980 12880
rect 21160 12680 23360 12880
rect 20980 12670 21160 12680
rect 18740 12400 18820 12410
rect 21260 12400 21340 12410
rect 16680 12160 18740 12400
rect 18820 12160 21260 12400
rect 18740 12150 18820 12160
rect 21260 12150 21340 12160
rect 17300 11940 17400 11950
rect 17480 11940 17560 11950
rect 20000 11940 20080 11950
rect 22520 11940 22600 11950
rect 16680 11820 17000 11830
rect 17400 11700 17480 11940
rect 17560 11700 20000 11940
rect 20080 11700 22520 11940
rect 22600 11700 22640 11940
rect 17300 11690 17400 11700
rect 17480 11690 17560 11700
rect 20000 11690 20080 11700
rect 16680 11670 17000 11680
rect 22240 10540 22640 11700
rect 22240 10160 25400 10540
rect 25060 9580 25400 10160
rect 25360 9180 25400 9580
rect 25360 9160 25380 9180
rect 25060 9150 25360 9160
<< via2 >>
rect 16680 13480 17000 13620
rect 20920 13100 21120 13360
rect 22840 13180 23100 13360
rect 16680 11680 17000 11820
<< metal3 >>
rect 16670 13620 17010 13625
rect 16670 13480 16680 13620
rect 17000 13480 17010 13620
rect 16670 13475 17010 13480
rect 16680 11825 17000 13475
rect 20910 13360 21130 13365
rect 22830 13360 23110 13365
rect 20910 13100 20920 13360
rect 21120 13180 22840 13360
rect 23100 13180 23120 13360
rect 21120 13100 23120 13180
rect 20910 13095 21130 13100
rect 16670 11820 17010 11825
rect 16670 11680 16680 11820
rect 17000 11680 17010 11820
rect 16670 11675 17010 11680
use isource_cmirror  isource_cmirror_0
timestamp 1645630008
transform 1 0 23200 0 1 12240
box 0 0 2044 2280
use isource_conv_tsmal  isource_conv_tsmal_0
timestamp 1645614240
transform 1 0 16700 0 1 6440
box 4250 6510 5820 8748
use isource_ref_transistor  isource_ref_transistor_0
timestamp 1645630008
transform 1 0 4813 0 1 12757
box -493 -117 12421 1103
use isource_ref_transistor  isource_ref_transistor_1
timestamp 1645630008
transform 1 0 4813 0 1 11547
box -493 -117 12421 1103
use sky130_fd_pr__nfet_01v8_834VMG  sky130_fd_pr__nfet_01v8_834VMG_0
timestamp 1645614240
transform 1 0 20043 0 1 12050
box -2683 -610 2683 610
use sky130_fd_pr__res_xhigh_po_1p41_JAGHGM  sky130_fd_pr__res_xhigh_po_1p41_JAGHGM_0
timestamp 1645614240
transform 1 0 24147 0 1 10578
box -1367 -1598 1367 1598
<< end >>
