magic
tech sky130A
magscale 1 2
timestamp 1647254192
<< error_p >>
rect -78 281 -20 287
rect 118 281 176 287
rect -78 247 -66 281
rect 118 247 130 281
rect -78 241 -20 247
rect 118 241 176 247
rect -176 -247 -118 -241
rect 20 -247 78 -241
rect -176 -281 -164 -247
rect 20 -281 32 -247
rect -176 -287 -118 -281
rect 20 -287 78 -281
<< nwell >>
rect -363 -419 363 419
<< pmos >>
rect -167 -200 -127 200
rect -69 -200 -29 200
rect 29 -200 69 200
rect 127 -200 167 200
<< pdiff >>
rect -225 188 -167 200
rect -225 -188 -213 188
rect -179 -188 -167 188
rect -225 -200 -167 -188
rect -127 188 -69 200
rect -127 -188 -115 188
rect -81 -188 -69 188
rect -127 -200 -69 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 69 188 127 200
rect 69 -188 81 188
rect 115 -188 127 188
rect 69 -200 127 -188
rect 167 188 225 200
rect 167 -188 179 188
rect 213 -188 225 188
rect 167 -200 225 -188
<< pdiffc >>
rect -213 -188 -179 188
rect -115 -188 -81 188
rect -17 -188 17 188
rect 81 -188 115 188
rect 179 -188 213 188
<< nsubdiff >>
rect -327 349 -231 383
rect 231 349 327 383
rect -327 287 -293 349
rect 293 287 327 349
rect -327 -349 -293 -287
rect 293 -349 327 -287
rect -327 -383 -231 -349
rect 231 -383 327 -349
<< nsubdiffcont >>
rect -231 349 231 383
rect -327 -287 -293 287
rect 293 -287 327 287
rect -231 -383 231 -349
<< poly >>
rect -82 281 -16 297
rect -82 247 -66 281
rect -32 247 -16 281
rect -82 231 -16 247
rect 114 281 180 297
rect 114 247 130 281
rect 164 247 180 281
rect 114 231 180 247
rect -167 200 -127 226
rect -69 200 -29 231
rect 29 200 69 226
rect 127 200 167 231
rect -167 -231 -127 -200
rect -69 -226 -29 -200
rect 29 -231 69 -200
rect 127 -226 167 -200
rect -180 -247 -114 -231
rect -180 -281 -164 -247
rect -130 -281 -114 -247
rect -180 -297 -114 -281
rect 16 -247 82 -231
rect 16 -281 32 -247
rect 66 -281 82 -247
rect 16 -297 82 -281
<< polycont >>
rect -66 247 -32 281
rect 130 247 164 281
rect -164 -281 -130 -247
rect 32 -281 66 -247
<< locali >>
rect -327 349 -231 383
rect 231 349 327 383
rect -327 287 -293 349
rect 293 287 327 349
rect -82 247 -66 281
rect -32 247 -16 281
rect 114 247 130 281
rect 164 247 180 281
rect -213 188 -179 204
rect -213 -204 -179 -188
rect -115 188 -81 204
rect -115 -204 -81 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 81 188 115 204
rect 81 -204 115 -188
rect 179 188 213 204
rect 179 -204 213 -188
rect -180 -281 -164 -247
rect -130 -281 -114 -247
rect 16 -281 32 -247
rect 66 -281 82 -247
rect -327 -349 -293 -287
rect 293 -349 327 -287
rect -327 -383 -231 -349
rect 231 -383 327 -349
<< viali >>
rect -66 247 -32 281
rect 130 247 164 281
rect -213 -188 -179 188
rect -115 -188 -81 188
rect -17 -188 17 188
rect 81 -188 115 188
rect 179 -188 213 188
rect -164 -281 -130 -247
rect 32 -281 66 -247
<< metal1 >>
rect -78 281 -20 287
rect -78 247 -66 281
rect -32 247 -20 281
rect -78 241 -20 247
rect 118 281 176 287
rect 118 247 130 281
rect 164 247 176 281
rect 118 241 176 247
rect -219 188 -173 200
rect -219 -188 -213 188
rect -179 -188 -173 188
rect -219 -200 -173 -188
rect -121 188 -75 200
rect -121 -188 -115 188
rect -81 -188 -75 188
rect -121 -200 -75 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 75 188 121 200
rect 75 -188 81 188
rect 115 -188 121 188
rect 75 -200 121 -188
rect 173 188 219 200
rect 173 -188 179 188
rect 213 -188 219 188
rect 173 -200 219 -188
rect -176 -247 -118 -241
rect -176 -281 -164 -247
rect -130 -281 -118 -247
rect -176 -287 -118 -281
rect 20 -247 78 -241
rect 20 -281 32 -247
rect 66 -281 78 -247
rect 20 -287 78 -281
<< properties >>
string FIXED_BBOX -310 -366 310 366
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 0.2 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
