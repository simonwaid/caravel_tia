magic
tech sky130A
magscale 1 2
timestamp 1646921651
<< pwell >>
rect -6457 -610 6457 610
<< nmos >>
rect -6261 -400 -5061 400
rect -5003 -400 -3803 400
rect -3745 -400 -2545 400
rect -2487 -400 -1287 400
rect -1229 -400 -29 400
rect 29 -400 1229 400
rect 1287 -400 2487 400
rect 2545 -400 3745 400
rect 3803 -400 5003 400
rect 5061 -400 6261 400
<< ndiff >>
rect -6319 388 -6261 400
rect -6319 -388 -6307 388
rect -6273 -388 -6261 388
rect -6319 -400 -6261 -388
rect -5061 388 -5003 400
rect -5061 -388 -5049 388
rect -5015 -388 -5003 388
rect -5061 -400 -5003 -388
rect -3803 388 -3745 400
rect -3803 -388 -3791 388
rect -3757 -388 -3745 388
rect -3803 -400 -3745 -388
rect -2545 388 -2487 400
rect -2545 -388 -2533 388
rect -2499 -388 -2487 388
rect -2545 -400 -2487 -388
rect -1287 388 -1229 400
rect -1287 -388 -1275 388
rect -1241 -388 -1229 388
rect -1287 -400 -1229 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 1229 388 1287 400
rect 1229 -388 1241 388
rect 1275 -388 1287 388
rect 1229 -400 1287 -388
rect 2487 388 2545 400
rect 2487 -388 2499 388
rect 2533 -388 2545 388
rect 2487 -400 2545 -388
rect 3745 388 3803 400
rect 3745 -388 3757 388
rect 3791 -388 3803 388
rect 3745 -400 3803 -388
rect 5003 388 5061 400
rect 5003 -388 5015 388
rect 5049 -388 5061 388
rect 5003 -400 5061 -388
rect 6261 388 6319 400
rect 6261 -388 6273 388
rect 6307 -388 6319 388
rect 6261 -400 6319 -388
<< ndiffc >>
rect -6307 -388 -6273 388
rect -5049 -388 -5015 388
rect -3791 -388 -3757 388
rect -2533 -388 -2499 388
rect -1275 -388 -1241 388
rect -17 -388 17 388
rect 1241 -388 1275 388
rect 2499 -388 2533 388
rect 3757 -388 3791 388
rect 5015 -388 5049 388
rect 6273 -388 6307 388
<< psubdiff >>
rect -6421 540 -6325 574
rect 6325 540 6421 574
rect -6421 478 -6387 540
rect 6387 478 6421 540
rect -6421 -540 -6387 -478
rect 6387 -540 6421 -478
rect -6421 -574 -6325 -540
rect 6325 -574 6421 -540
<< psubdiffcont >>
rect -6325 540 6325 574
rect -6421 -478 -6387 478
rect 6387 -478 6421 478
rect -6325 -574 6325 -540
<< poly >>
rect -6261 472 -5061 488
rect -6261 438 -6245 472
rect -5077 438 -5061 472
rect -6261 400 -5061 438
rect -5003 472 -3803 488
rect -5003 438 -4987 472
rect -3819 438 -3803 472
rect -5003 400 -3803 438
rect -3745 472 -2545 488
rect -3745 438 -3729 472
rect -2561 438 -2545 472
rect -3745 400 -2545 438
rect -2487 472 -1287 488
rect -2487 438 -2471 472
rect -1303 438 -1287 472
rect -2487 400 -1287 438
rect -1229 472 -29 488
rect -1229 438 -1213 472
rect -45 438 -29 472
rect -1229 400 -29 438
rect 29 472 1229 488
rect 29 438 45 472
rect 1213 438 1229 472
rect 29 400 1229 438
rect 1287 472 2487 488
rect 1287 438 1303 472
rect 2471 438 2487 472
rect 1287 400 2487 438
rect 2545 472 3745 488
rect 2545 438 2561 472
rect 3729 438 3745 472
rect 2545 400 3745 438
rect 3803 472 5003 488
rect 3803 438 3819 472
rect 4987 438 5003 472
rect 3803 400 5003 438
rect 5061 472 6261 488
rect 5061 438 5077 472
rect 6245 438 6261 472
rect 5061 400 6261 438
rect -6261 -438 -5061 -400
rect -6261 -472 -6245 -438
rect -5077 -472 -5061 -438
rect -6261 -488 -5061 -472
rect -5003 -438 -3803 -400
rect -5003 -472 -4987 -438
rect -3819 -472 -3803 -438
rect -5003 -488 -3803 -472
rect -3745 -438 -2545 -400
rect -3745 -472 -3729 -438
rect -2561 -472 -2545 -438
rect -3745 -488 -2545 -472
rect -2487 -438 -1287 -400
rect -2487 -472 -2471 -438
rect -1303 -472 -1287 -438
rect -2487 -488 -1287 -472
rect -1229 -438 -29 -400
rect -1229 -472 -1213 -438
rect -45 -472 -29 -438
rect -1229 -488 -29 -472
rect 29 -438 1229 -400
rect 29 -472 45 -438
rect 1213 -472 1229 -438
rect 29 -488 1229 -472
rect 1287 -438 2487 -400
rect 1287 -472 1303 -438
rect 2471 -472 2487 -438
rect 1287 -488 2487 -472
rect 2545 -438 3745 -400
rect 2545 -472 2561 -438
rect 3729 -472 3745 -438
rect 2545 -488 3745 -472
rect 3803 -438 5003 -400
rect 3803 -472 3819 -438
rect 4987 -472 5003 -438
rect 3803 -488 5003 -472
rect 5061 -438 6261 -400
rect 5061 -472 5077 -438
rect 6245 -472 6261 -438
rect 5061 -488 6261 -472
<< polycont >>
rect -6245 438 -5077 472
rect -4987 438 -3819 472
rect -3729 438 -2561 472
rect -2471 438 -1303 472
rect -1213 438 -45 472
rect 45 438 1213 472
rect 1303 438 2471 472
rect 2561 438 3729 472
rect 3819 438 4987 472
rect 5077 438 6245 472
rect -6245 -472 -5077 -438
rect -4987 -472 -3819 -438
rect -3729 -472 -2561 -438
rect -2471 -472 -1303 -438
rect -1213 -472 -45 -438
rect 45 -472 1213 -438
rect 1303 -472 2471 -438
rect 2561 -472 3729 -438
rect 3819 -472 4987 -438
rect 5077 -472 6245 -438
<< locali >>
rect -6421 540 -6325 574
rect 6325 540 6421 574
rect -6421 478 -6387 540
rect 6387 478 6421 540
rect -6261 438 -6245 472
rect -5077 438 -5061 472
rect -5003 438 -4987 472
rect -3819 438 -3803 472
rect -3745 438 -3729 472
rect -2561 438 -2545 472
rect -2487 438 -2471 472
rect -1303 438 -1287 472
rect -1229 438 -1213 472
rect -45 438 -29 472
rect 29 438 45 472
rect 1213 438 1229 472
rect 1287 438 1303 472
rect 2471 438 2487 472
rect 2545 438 2561 472
rect 3729 438 3745 472
rect 3803 438 3819 472
rect 4987 438 5003 472
rect 5061 438 5077 472
rect 6245 438 6261 472
rect -6307 388 -6273 404
rect -6307 -404 -6273 -388
rect -5049 388 -5015 404
rect -5049 -404 -5015 -388
rect -3791 388 -3757 404
rect -3791 -404 -3757 -388
rect -2533 388 -2499 404
rect -2533 -404 -2499 -388
rect -1275 388 -1241 404
rect -1275 -404 -1241 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 1241 388 1275 404
rect 1241 -404 1275 -388
rect 2499 388 2533 404
rect 2499 -404 2533 -388
rect 3757 388 3791 404
rect 3757 -404 3791 -388
rect 5015 388 5049 404
rect 5015 -404 5049 -388
rect 6273 388 6307 404
rect 6273 -404 6307 -388
rect -6261 -472 -6245 -438
rect -5077 -472 -5061 -438
rect -5003 -472 -4987 -438
rect -3819 -472 -3803 -438
rect -3745 -472 -3729 -438
rect -2561 -472 -2545 -438
rect -2487 -472 -2471 -438
rect -1303 -472 -1287 -438
rect -1229 -472 -1213 -438
rect -45 -472 -29 -438
rect 29 -472 45 -438
rect 1213 -472 1229 -438
rect 1287 -472 1303 -438
rect 2471 -472 2487 -438
rect 2545 -472 2561 -438
rect 3729 -472 3745 -438
rect 3803 -472 3819 -438
rect 4987 -472 5003 -438
rect 5061 -472 5077 -438
rect 6245 -472 6261 -438
rect -6421 -540 -6387 -478
rect 6387 -540 6421 -478
rect -6421 -574 -6325 -540
rect 6325 -574 6421 -540
<< viali >>
rect -6245 438 -5077 472
rect -4987 438 -3819 472
rect -3729 438 -2561 472
rect -2471 438 -1303 472
rect -1213 438 -45 472
rect 45 438 1213 472
rect 1303 438 2471 472
rect 2561 438 3729 472
rect 3819 438 4987 472
rect 5077 438 6245 472
rect -6307 -388 -6273 388
rect -5049 -388 -5015 388
rect -3791 -388 -3757 388
rect -2533 -388 -2499 388
rect -1275 -388 -1241 388
rect -17 -388 17 388
rect 1241 -388 1275 388
rect 2499 -388 2533 388
rect 3757 -388 3791 388
rect 5015 -388 5049 388
rect 6273 -388 6307 388
rect -6245 -472 -5077 -438
rect -4987 -472 -3819 -438
rect -3729 -472 -2561 -438
rect -2471 -472 -1303 -438
rect -1213 -472 -45 -438
rect 45 -472 1213 -438
rect 1303 -472 2471 -438
rect 2561 -472 3729 -438
rect 3819 -472 4987 -438
rect 5077 -472 6245 -438
<< metal1 >>
rect -6257 472 -5065 478
rect -6257 438 -6245 472
rect -5077 438 -5065 472
rect -6257 432 -5065 438
rect -4999 472 -3807 478
rect -4999 438 -4987 472
rect -3819 438 -3807 472
rect -4999 432 -3807 438
rect -3741 472 -2549 478
rect -3741 438 -3729 472
rect -2561 438 -2549 472
rect -3741 432 -2549 438
rect -2483 472 -1291 478
rect -2483 438 -2471 472
rect -1303 438 -1291 472
rect -2483 432 -1291 438
rect -1225 472 -33 478
rect -1225 438 -1213 472
rect -45 438 -33 472
rect -1225 432 -33 438
rect 33 472 1225 478
rect 33 438 45 472
rect 1213 438 1225 472
rect 33 432 1225 438
rect 1291 472 2483 478
rect 1291 438 1303 472
rect 2471 438 2483 472
rect 1291 432 2483 438
rect 2549 472 3741 478
rect 2549 438 2561 472
rect 3729 438 3741 472
rect 2549 432 3741 438
rect 3807 472 4999 478
rect 3807 438 3819 472
rect 4987 438 4999 472
rect 3807 432 4999 438
rect 5065 472 6257 478
rect 5065 438 5077 472
rect 6245 438 6257 472
rect 5065 432 6257 438
rect -6313 388 -6267 400
rect -6313 -388 -6307 388
rect -6273 -388 -6267 388
rect -6313 -400 -6267 -388
rect -5055 388 -5009 400
rect -5055 -388 -5049 388
rect -5015 -388 -5009 388
rect -5055 -400 -5009 -388
rect -3797 388 -3751 400
rect -3797 -388 -3791 388
rect -3757 -388 -3751 388
rect -3797 -400 -3751 -388
rect -2539 388 -2493 400
rect -2539 -388 -2533 388
rect -2499 -388 -2493 388
rect -2539 -400 -2493 -388
rect -1281 388 -1235 400
rect -1281 -388 -1275 388
rect -1241 -388 -1235 388
rect -1281 -400 -1235 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 1235 388 1281 400
rect 1235 -388 1241 388
rect 1275 -388 1281 388
rect 1235 -400 1281 -388
rect 2493 388 2539 400
rect 2493 -388 2499 388
rect 2533 -388 2539 388
rect 2493 -400 2539 -388
rect 3751 388 3797 400
rect 3751 -388 3757 388
rect 3791 -388 3797 388
rect 3751 -400 3797 -388
rect 5009 388 5055 400
rect 5009 -388 5015 388
rect 5049 -388 5055 388
rect 5009 -400 5055 -388
rect 6267 388 6313 400
rect 6267 -388 6273 388
rect 6307 -388 6313 388
rect 6267 -400 6313 -388
rect -6257 -438 -5065 -432
rect -6257 -472 -6245 -438
rect -5077 -472 -5065 -438
rect -6257 -478 -5065 -472
rect -4999 -438 -3807 -432
rect -4999 -472 -4987 -438
rect -3819 -472 -3807 -438
rect -4999 -478 -3807 -472
rect -3741 -438 -2549 -432
rect -3741 -472 -3729 -438
rect -2561 -472 -2549 -438
rect -3741 -478 -2549 -472
rect -2483 -438 -1291 -432
rect -2483 -472 -2471 -438
rect -1303 -472 -1291 -438
rect -2483 -478 -1291 -472
rect -1225 -438 -33 -432
rect -1225 -472 -1213 -438
rect -45 -472 -33 -438
rect -1225 -478 -33 -472
rect 33 -438 1225 -432
rect 33 -472 45 -438
rect 1213 -472 1225 -438
rect 33 -478 1225 -472
rect 1291 -438 2483 -432
rect 1291 -472 1303 -438
rect 2471 -472 2483 -438
rect 1291 -478 2483 -472
rect 2549 -438 3741 -432
rect 2549 -472 2561 -438
rect 3729 -472 3741 -438
rect 2549 -478 3741 -472
rect 3807 -438 4999 -432
rect 3807 -472 3819 -438
rect 4987 -472 4999 -438
rect 3807 -478 4999 -472
rect 5065 -438 6257 -432
rect 5065 -472 5077 -438
rect 6245 -472 6257 -438
rect 5065 -478 6257 -472
<< properties >>
string FIXED_BBOX -6404 -557 6404 557
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 4 l 6 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
