magic
tech sky130A
magscale 1 2
timestamp 1646921651
<< nwell >>
rect 623 1186 2061 1252
rect 2421 1186 3859 1252
rect 734 1180 774 1186
rect 930 1180 970 1186
rect 1126 1180 1166 1186
rect 1322 1180 1362 1186
rect 1518 1180 1558 1186
rect 1714 1180 1754 1186
rect 1910 1180 1950 1186
rect 2532 1180 2572 1186
rect 2728 1180 2768 1186
rect 2924 1180 2964 1186
rect 3120 1180 3160 1186
rect 3316 1180 3356 1186
rect 3512 1180 3552 1186
rect 3708 1180 3748 1186
rect 636 724 676 730
rect 832 724 872 730
rect 1028 724 1068 730
rect 1224 724 1264 730
rect 1420 724 1460 730
rect 1616 724 1656 730
rect 1812 724 1852 730
rect 2008 724 2048 730
rect 2434 724 2474 730
rect 2630 724 2670 730
rect 2826 724 2866 730
rect 3022 724 3062 730
rect 3218 724 3258 730
rect 3414 724 3454 730
rect 3610 724 3650 730
rect 3806 724 3846 730
rect 623 658 2061 724
rect 2421 658 3859 724
rect 623 550 2061 616
rect 2421 550 3859 616
rect 636 544 676 550
rect 832 544 872 550
rect 1028 544 1068 550
rect 1224 544 1264 550
rect 1420 544 1460 550
rect 1616 544 1656 550
rect 1812 544 1852 550
rect 2008 544 2048 550
rect 2434 544 2474 550
rect 2630 544 2670 550
rect 2826 544 2866 550
rect 3022 544 3062 550
rect 3218 544 3258 550
rect 3414 544 3454 550
rect 3610 544 3650 550
rect 3806 544 3846 550
rect 734 88 774 94
rect 930 88 970 94
rect 1126 88 1166 94
rect 1322 88 1362 94
rect 1518 88 1558 94
rect 1714 88 1754 94
rect 1910 88 1950 94
rect 2532 88 2572 94
rect 2728 88 2768 94
rect 2924 88 2964 94
rect 3120 88 3160 94
rect 3316 88 3356 94
rect 3512 88 3552 94
rect 3708 88 3748 94
rect 623 22 2061 88
rect 2421 22 3859 88
<< poly >>
rect 623 1236 2061 1252
rect 623 1202 737 1236
rect 771 1202 933 1236
rect 967 1202 1129 1236
rect 1163 1202 1325 1236
rect 1359 1202 1521 1236
rect 1555 1202 1717 1236
rect 1751 1202 1913 1236
rect 1947 1202 2061 1236
rect 623 1186 2061 1202
rect 2421 1236 3859 1252
rect 2421 1202 2535 1236
rect 2569 1202 2731 1236
rect 2765 1202 2927 1236
rect 2961 1202 3123 1236
rect 3157 1202 3319 1236
rect 3353 1202 3515 1236
rect 3549 1202 3711 1236
rect 3745 1202 3859 1236
rect 2421 1186 3859 1202
rect 734 1180 774 1186
rect 930 1180 970 1186
rect 1126 1180 1166 1186
rect 1322 1180 1362 1186
rect 1518 1180 1558 1186
rect 1714 1180 1754 1186
rect 1910 1180 1950 1186
rect 2532 1180 2572 1186
rect 2728 1180 2768 1186
rect 2924 1180 2964 1186
rect 3120 1180 3160 1186
rect 3316 1180 3356 1186
rect 3512 1180 3552 1186
rect 3708 1180 3748 1186
rect 636 724 676 730
rect 832 724 872 730
rect 1028 724 1068 730
rect 1224 724 1264 730
rect 1420 724 1460 730
rect 1616 724 1656 730
rect 1812 724 1852 730
rect 2008 724 2048 730
rect 2434 724 2474 730
rect 2630 724 2670 730
rect 2826 724 2866 730
rect 3022 724 3062 730
rect 3218 724 3258 730
rect 3414 724 3454 730
rect 3610 724 3650 730
rect 3806 724 3846 730
rect 623 708 2061 724
rect 623 674 639 708
rect 673 674 835 708
rect 869 674 1031 708
rect 1065 674 1227 708
rect 1261 674 1423 708
rect 1457 674 1619 708
rect 1653 674 1815 708
rect 1849 674 2011 708
rect 2045 674 2061 708
rect 623 658 2061 674
rect 2421 708 3859 724
rect 2421 674 2437 708
rect 2471 674 2633 708
rect 2667 674 2829 708
rect 2863 674 3025 708
rect 3059 674 3221 708
rect 3255 674 3417 708
rect 3451 674 3613 708
rect 3647 674 3809 708
rect 3843 674 3859 708
rect 2421 658 3859 674
rect 623 600 2061 616
rect 623 566 639 600
rect 673 566 835 600
rect 869 566 1031 600
rect 1065 566 1227 600
rect 1261 566 1423 600
rect 1457 566 1619 600
rect 1653 566 1815 600
rect 1849 566 2011 600
rect 2045 566 2061 600
rect 623 550 2061 566
rect 2421 600 3859 616
rect 2421 566 2437 600
rect 2471 566 2633 600
rect 2667 566 2829 600
rect 2863 566 3025 600
rect 3059 566 3221 600
rect 3255 566 3417 600
rect 3451 566 3613 600
rect 3647 566 3809 600
rect 3843 566 3859 600
rect 2421 550 3859 566
rect 636 544 676 550
rect 832 544 872 550
rect 1028 544 1068 550
rect 1224 544 1264 550
rect 1420 544 1460 550
rect 1616 544 1656 550
rect 1812 544 1852 550
rect 2008 544 2048 550
rect 2434 544 2474 550
rect 2630 544 2670 550
rect 2826 544 2866 550
rect 3022 544 3062 550
rect 3218 544 3258 550
rect 3414 544 3454 550
rect 3610 544 3650 550
rect 3806 544 3846 550
rect 734 88 774 94
rect 930 88 970 94
rect 1126 88 1166 94
rect 1322 88 1362 94
rect 1518 88 1558 94
rect 1714 88 1754 94
rect 1910 88 1950 94
rect 2532 88 2572 94
rect 2728 88 2768 94
rect 2924 88 2964 94
rect 3120 88 3160 94
rect 3316 88 3356 94
rect 3512 88 3552 94
rect 3708 88 3748 94
rect 623 72 2061 88
rect 623 38 737 72
rect 771 38 933 72
rect 967 38 1129 72
rect 1163 38 1325 72
rect 1359 38 1521 72
rect 1555 38 1717 72
rect 1751 38 1913 72
rect 1947 38 2061 72
rect 623 22 2061 38
rect 2421 72 3859 88
rect 2421 38 2535 72
rect 2569 38 2731 72
rect 2765 38 2927 72
rect 2961 38 3123 72
rect 3157 38 3319 72
rect 3353 38 3515 72
rect 3549 38 3711 72
rect 3745 38 3859 72
rect 2421 22 3859 38
rect 622 -240 3040 -224
rect 622 -274 736 -240
rect 770 -274 932 -240
rect 966 -274 1128 -240
rect 1162 -274 1324 -240
rect 1358 -274 1520 -240
rect 1554 -274 1716 -240
rect 1750 -274 1912 -240
rect 1946 -274 2108 -240
rect 2142 -274 2304 -240
rect 2338 -274 2500 -240
rect 2534 -274 2696 -240
rect 2730 -274 2892 -240
rect 2926 -274 3040 -240
rect 622 -290 3040 -274
rect 622 -750 3040 -734
rect 622 -784 638 -750
rect 672 -784 834 -750
rect 868 -784 1030 -750
rect 1064 -784 1226 -750
rect 1260 -784 1422 -750
rect 1456 -784 1618 -750
rect 1652 -784 1814 -750
rect 1848 -784 2010 -750
rect 2044 -784 2206 -750
rect 2240 -784 2402 -750
rect 2436 -784 2598 -750
rect 2632 -784 2794 -750
rect 2828 -784 2990 -750
rect 3024 -784 3040 -750
rect 622 -800 3040 -784
rect 623 -858 3041 -842
rect 623 -892 639 -858
rect 673 -892 835 -858
rect 869 -892 1031 -858
rect 1065 -892 1227 -858
rect 1261 -892 1423 -858
rect 1457 -892 1619 -858
rect 1653 -892 1815 -858
rect 1849 -892 2011 -858
rect 2045 -892 2207 -858
rect 2241 -892 2403 -858
rect 2437 -892 2599 -858
rect 2633 -892 2795 -858
rect 2829 -892 2991 -858
rect 3025 -892 3041 -858
rect 623 -908 3041 -892
rect 623 -1368 3041 -1352
rect 623 -1402 737 -1368
rect 771 -1402 933 -1368
rect 967 -1402 1129 -1368
rect 1163 -1402 1325 -1368
rect 1359 -1402 1521 -1368
rect 1555 -1402 1717 -1368
rect 1751 -1402 1913 -1368
rect 1947 -1402 2109 -1368
rect 2143 -1402 2305 -1368
rect 2339 -1402 2501 -1368
rect 2535 -1402 2697 -1368
rect 2731 -1402 2893 -1368
rect 2927 -1402 3041 -1368
rect 623 -1418 3041 -1402
rect 622 -1684 3040 -1668
rect 622 -1718 736 -1684
rect 770 -1718 932 -1684
rect 966 -1718 1128 -1684
rect 1162 -1718 1324 -1684
rect 1358 -1718 1520 -1684
rect 1554 -1718 1716 -1684
rect 1750 -1718 1912 -1684
rect 1946 -1718 2108 -1684
rect 2142 -1718 2304 -1684
rect 2338 -1718 2500 -1684
rect 2534 -1718 2696 -1684
rect 2730 -1718 2892 -1684
rect 2926 -1718 3040 -1684
rect 622 -1734 3040 -1718
rect 622 -2194 3040 -2178
rect 622 -2228 638 -2194
rect 672 -2228 834 -2194
rect 868 -2228 1030 -2194
rect 1064 -2228 1226 -2194
rect 1260 -2228 1422 -2194
rect 1456 -2228 1618 -2194
rect 1652 -2228 1814 -2194
rect 1848 -2228 2010 -2194
rect 2044 -2228 2206 -2194
rect 2240 -2228 2402 -2194
rect 2436 -2228 2598 -2194
rect 2632 -2228 2794 -2194
rect 2828 -2228 2990 -2194
rect 3024 -2228 3040 -2194
rect 622 -2244 3040 -2228
rect 623 -2302 3041 -2286
rect 623 -2336 639 -2302
rect 673 -2336 835 -2302
rect 869 -2336 1031 -2302
rect 1065 -2336 1227 -2302
rect 1261 -2336 1423 -2302
rect 1457 -2336 1619 -2302
rect 1653 -2336 1815 -2302
rect 1849 -2336 2011 -2302
rect 2045 -2336 2207 -2302
rect 2241 -2336 2403 -2302
rect 2437 -2336 2599 -2302
rect 2633 -2336 2795 -2302
rect 2829 -2336 2991 -2302
rect 3025 -2336 3041 -2302
rect 623 -2352 3041 -2336
rect 623 -2812 3041 -2796
rect 623 -2846 737 -2812
rect 771 -2846 933 -2812
rect 967 -2846 1129 -2812
rect 1163 -2846 1325 -2812
rect 1359 -2846 1521 -2812
rect 1555 -2846 1717 -2812
rect 1751 -2846 1913 -2812
rect 1947 -2846 2109 -2812
rect 2143 -2846 2305 -2812
rect 2339 -2846 2501 -2812
rect 2535 -2846 2697 -2812
rect 2731 -2846 2893 -2812
rect 2927 -2846 3041 -2812
rect 623 -2862 3041 -2846
<< polycont >>
rect 737 1202 771 1236
rect 933 1202 967 1236
rect 1129 1202 1163 1236
rect 1325 1202 1359 1236
rect 1521 1202 1555 1236
rect 1717 1202 1751 1236
rect 1913 1202 1947 1236
rect 2535 1202 2569 1236
rect 2731 1202 2765 1236
rect 2927 1202 2961 1236
rect 3123 1202 3157 1236
rect 3319 1202 3353 1236
rect 3515 1202 3549 1236
rect 3711 1202 3745 1236
rect 639 674 673 708
rect 835 674 869 708
rect 1031 674 1065 708
rect 1227 674 1261 708
rect 1423 674 1457 708
rect 1619 674 1653 708
rect 1815 674 1849 708
rect 2011 674 2045 708
rect 2437 674 2471 708
rect 2633 674 2667 708
rect 2829 674 2863 708
rect 3025 674 3059 708
rect 3221 674 3255 708
rect 3417 674 3451 708
rect 3613 674 3647 708
rect 3809 674 3843 708
rect 639 566 673 600
rect 835 566 869 600
rect 1031 566 1065 600
rect 1227 566 1261 600
rect 1423 566 1457 600
rect 1619 566 1653 600
rect 1815 566 1849 600
rect 2011 566 2045 600
rect 2437 566 2471 600
rect 2633 566 2667 600
rect 2829 566 2863 600
rect 3025 566 3059 600
rect 3221 566 3255 600
rect 3417 566 3451 600
rect 3613 566 3647 600
rect 3809 566 3843 600
rect 737 38 771 72
rect 933 38 967 72
rect 1129 38 1163 72
rect 1325 38 1359 72
rect 1521 38 1555 72
rect 1717 38 1751 72
rect 1913 38 1947 72
rect 2535 38 2569 72
rect 2731 38 2765 72
rect 2927 38 2961 72
rect 3123 38 3157 72
rect 3319 38 3353 72
rect 3515 38 3549 72
rect 3711 38 3745 72
rect 736 -274 770 -240
rect 932 -274 966 -240
rect 1128 -274 1162 -240
rect 1324 -274 1358 -240
rect 1520 -274 1554 -240
rect 1716 -274 1750 -240
rect 1912 -274 1946 -240
rect 2108 -274 2142 -240
rect 2304 -274 2338 -240
rect 2500 -274 2534 -240
rect 2696 -274 2730 -240
rect 2892 -274 2926 -240
rect 638 -784 672 -750
rect 834 -784 868 -750
rect 1030 -784 1064 -750
rect 1226 -784 1260 -750
rect 1422 -784 1456 -750
rect 1618 -784 1652 -750
rect 1814 -784 1848 -750
rect 2010 -784 2044 -750
rect 2206 -784 2240 -750
rect 2402 -784 2436 -750
rect 2598 -784 2632 -750
rect 2794 -784 2828 -750
rect 2990 -784 3024 -750
rect 639 -892 673 -858
rect 835 -892 869 -858
rect 1031 -892 1065 -858
rect 1227 -892 1261 -858
rect 1423 -892 1457 -858
rect 1619 -892 1653 -858
rect 1815 -892 1849 -858
rect 2011 -892 2045 -858
rect 2207 -892 2241 -858
rect 2403 -892 2437 -858
rect 2599 -892 2633 -858
rect 2795 -892 2829 -858
rect 2991 -892 3025 -858
rect 737 -1402 771 -1368
rect 933 -1402 967 -1368
rect 1129 -1402 1163 -1368
rect 1325 -1402 1359 -1368
rect 1521 -1402 1555 -1368
rect 1717 -1402 1751 -1368
rect 1913 -1402 1947 -1368
rect 2109 -1402 2143 -1368
rect 2305 -1402 2339 -1368
rect 2501 -1402 2535 -1368
rect 2697 -1402 2731 -1368
rect 2893 -1402 2927 -1368
rect 736 -1718 770 -1684
rect 932 -1718 966 -1684
rect 1128 -1718 1162 -1684
rect 1324 -1718 1358 -1684
rect 1520 -1718 1554 -1684
rect 1716 -1718 1750 -1684
rect 1912 -1718 1946 -1684
rect 2108 -1718 2142 -1684
rect 2304 -1718 2338 -1684
rect 2500 -1718 2534 -1684
rect 2696 -1718 2730 -1684
rect 2892 -1718 2926 -1684
rect 638 -2228 672 -2194
rect 834 -2228 868 -2194
rect 1030 -2228 1064 -2194
rect 1226 -2228 1260 -2194
rect 1422 -2228 1456 -2194
rect 1618 -2228 1652 -2194
rect 1814 -2228 1848 -2194
rect 2010 -2228 2044 -2194
rect 2206 -2228 2240 -2194
rect 2402 -2228 2436 -2194
rect 2598 -2228 2632 -2194
rect 2794 -2228 2828 -2194
rect 2990 -2228 3024 -2194
rect 639 -2336 673 -2302
rect 835 -2336 869 -2302
rect 1031 -2336 1065 -2302
rect 1227 -2336 1261 -2302
rect 1423 -2336 1457 -2302
rect 1619 -2336 1653 -2302
rect 1815 -2336 1849 -2302
rect 2011 -2336 2045 -2302
rect 2207 -2336 2241 -2302
rect 2403 -2336 2437 -2302
rect 2599 -2336 2633 -2302
rect 2795 -2336 2829 -2302
rect 2991 -2336 3025 -2302
rect 737 -2846 771 -2812
rect 933 -2846 967 -2812
rect 1129 -2846 1163 -2812
rect 1325 -2846 1359 -2812
rect 1521 -2846 1555 -2812
rect 1717 -2846 1751 -2812
rect 1913 -2846 1947 -2812
rect 2109 -2846 2143 -2812
rect 2305 -2846 2339 -2812
rect 2501 -2846 2535 -2812
rect 2697 -2846 2731 -2812
rect 2893 -2846 2927 -2812
<< locali >>
rect 623 1202 737 1236
rect 771 1202 933 1236
rect 967 1202 1129 1236
rect 1163 1202 1325 1236
rect 1359 1202 1521 1236
rect 1555 1202 1717 1236
rect 1751 1202 1913 1236
rect 1947 1202 2061 1236
rect 2421 1202 2535 1236
rect 2569 1202 2731 1236
rect 2765 1202 2927 1236
rect 2961 1202 3123 1236
rect 3157 1202 3319 1236
rect 3353 1202 3515 1236
rect 3549 1202 3711 1236
rect 3745 1202 3859 1236
rect 623 674 639 708
rect 673 674 835 708
rect 869 674 1031 708
rect 1065 674 1227 708
rect 1261 674 1423 708
rect 1457 674 1619 708
rect 1653 674 1815 708
rect 1849 674 2011 708
rect 2045 674 2061 708
rect 2421 674 2437 708
rect 2471 674 2633 708
rect 2667 674 2829 708
rect 2863 674 3025 708
rect 3059 674 3221 708
rect 3255 674 3417 708
rect 3451 674 3613 708
rect 3647 674 3809 708
rect 3843 674 3859 708
rect 623 566 639 600
rect 673 566 835 600
rect 869 566 1031 600
rect 1065 566 1227 600
rect 1261 566 1423 600
rect 1457 566 1619 600
rect 1653 566 1815 600
rect 1849 566 2011 600
rect 2045 566 2061 600
rect 2421 566 2437 600
rect 2471 566 2633 600
rect 2667 566 2829 600
rect 2863 566 3025 600
rect 3059 566 3221 600
rect 3255 566 3417 600
rect 3451 566 3613 600
rect 3647 566 3809 600
rect 3843 566 3859 600
rect 623 38 737 72
rect 771 38 933 72
rect 967 38 1129 72
rect 1163 38 1325 72
rect 1359 38 1521 72
rect 1555 38 1717 72
rect 1751 38 1913 72
rect 1947 38 2061 72
rect 2421 38 2535 72
rect 2569 38 2731 72
rect 2765 38 2927 72
rect 2961 38 3123 72
rect 3157 38 3319 72
rect 3353 38 3515 72
rect 3549 38 3711 72
rect 3745 38 3859 72
rect 622 -274 736 -240
rect 770 -274 932 -240
rect 966 -274 1128 -240
rect 1162 -274 1324 -240
rect 1358 -274 1520 -240
rect 1554 -274 1716 -240
rect 1750 -274 1912 -240
rect 1946 -274 2108 -240
rect 2142 -274 2304 -240
rect 2338 -274 2500 -240
rect 2534 -274 2696 -240
rect 2730 -274 2892 -240
rect 2926 -274 3040 -240
rect 622 -784 638 -750
rect 672 -784 834 -750
rect 868 -784 1030 -750
rect 1064 -784 1226 -750
rect 1260 -784 1422 -750
rect 1456 -784 1618 -750
rect 1652 -784 1814 -750
rect 1848 -784 2010 -750
rect 2044 -784 2206 -750
rect 2240 -784 2402 -750
rect 2436 -784 2598 -750
rect 2632 -784 2794 -750
rect 2828 -784 2990 -750
rect 3024 -784 3040 -750
rect 623 -892 639 -858
rect 673 -892 835 -858
rect 869 -892 1031 -858
rect 1065 -892 1227 -858
rect 1261 -892 1423 -858
rect 1457 -892 1619 -858
rect 1653 -892 1815 -858
rect 1849 -892 2011 -858
rect 2045 -892 2207 -858
rect 2241 -892 2403 -858
rect 2437 -892 2599 -858
rect 2633 -892 2795 -858
rect 2829 -892 2991 -858
rect 3025 -892 3041 -858
rect 623 -1402 737 -1368
rect 771 -1402 933 -1368
rect 967 -1402 1129 -1368
rect 1163 -1402 1325 -1368
rect 1359 -1402 1521 -1368
rect 1555 -1402 1717 -1368
rect 1751 -1402 1913 -1368
rect 1947 -1402 2109 -1368
rect 2143 -1402 2305 -1368
rect 2339 -1402 2501 -1368
rect 2535 -1402 2697 -1368
rect 2731 -1402 2893 -1368
rect 2927 -1402 3041 -1368
rect 622 -1718 736 -1684
rect 770 -1718 932 -1684
rect 966 -1718 1128 -1684
rect 1162 -1718 1324 -1684
rect 1358 -1718 1520 -1684
rect 1554 -1718 1716 -1684
rect 1750 -1718 1912 -1684
rect 1946 -1718 2108 -1684
rect 2142 -1718 2304 -1684
rect 2338 -1718 2500 -1684
rect 2534 -1718 2696 -1684
rect 2730 -1718 2892 -1684
rect 2926 -1718 3040 -1684
rect 622 -2228 638 -2194
rect 672 -2228 834 -2194
rect 868 -2228 1030 -2194
rect 1064 -2228 1226 -2194
rect 1260 -2228 1422 -2194
rect 1456 -2228 1618 -2194
rect 1652 -2228 1814 -2194
rect 1848 -2228 2010 -2194
rect 2044 -2228 2206 -2194
rect 2240 -2228 2402 -2194
rect 2436 -2228 2598 -2194
rect 2632 -2228 2794 -2194
rect 2828 -2228 2990 -2194
rect 3024 -2228 3040 -2194
rect 623 -2336 639 -2302
rect 673 -2336 835 -2302
rect 869 -2336 1031 -2302
rect 1065 -2336 1227 -2302
rect 1261 -2336 1423 -2302
rect 1457 -2336 1619 -2302
rect 1653 -2336 1815 -2302
rect 1849 -2336 2011 -2302
rect 2045 -2336 2207 -2302
rect 2241 -2336 2403 -2302
rect 2437 -2336 2599 -2302
rect 2633 -2336 2795 -2302
rect 2829 -2336 2991 -2302
rect 3025 -2336 3041 -2302
rect 623 -2846 737 -2812
rect 771 -2846 933 -2812
rect 967 -2846 1129 -2812
rect 1163 -2846 1325 -2812
rect 1359 -2846 1521 -2812
rect 1555 -2846 1717 -2812
rect 1751 -2846 1913 -2812
rect 1947 -2846 2109 -2812
rect 2143 -2846 2305 -2812
rect 2339 -2846 2501 -2812
rect 2535 -2846 2697 -2812
rect 2731 -2846 2893 -2812
rect 2927 -2846 3041 -2812
<< viali >>
rect 737 1202 771 1236
rect 933 1202 967 1236
rect 1129 1202 1163 1236
rect 1325 1202 1359 1236
rect 1521 1202 1555 1236
rect 1717 1202 1751 1236
rect 1913 1202 1947 1236
rect 2535 1202 2569 1236
rect 2731 1202 2765 1236
rect 2927 1202 2961 1236
rect 3123 1202 3157 1236
rect 3319 1202 3353 1236
rect 3515 1202 3549 1236
rect 3711 1202 3745 1236
rect 639 674 673 708
rect 835 674 869 708
rect 1031 674 1065 708
rect 1227 674 1261 708
rect 1423 674 1457 708
rect 1619 674 1653 708
rect 1815 674 1849 708
rect 2011 674 2045 708
rect 2437 674 2471 708
rect 2633 674 2667 708
rect 2829 674 2863 708
rect 3025 674 3059 708
rect 3221 674 3255 708
rect 3417 674 3451 708
rect 3613 674 3647 708
rect 3809 674 3843 708
rect 639 566 673 600
rect 835 566 869 600
rect 1031 566 1065 600
rect 1227 566 1261 600
rect 1423 566 1457 600
rect 1619 566 1653 600
rect 1815 566 1849 600
rect 2011 566 2045 600
rect 2437 566 2471 600
rect 2633 566 2667 600
rect 2829 566 2863 600
rect 3025 566 3059 600
rect 3221 566 3255 600
rect 3417 566 3451 600
rect 3613 566 3647 600
rect 3809 566 3843 600
rect 737 38 771 72
rect 933 38 967 72
rect 1129 38 1163 72
rect 1325 38 1359 72
rect 1521 38 1555 72
rect 1717 38 1751 72
rect 1913 38 1947 72
rect 2535 38 2569 72
rect 2731 38 2765 72
rect 2927 38 2961 72
rect 3123 38 3157 72
rect 3319 38 3353 72
rect 3515 38 3549 72
rect 3711 38 3745 72
rect 736 -274 770 -240
rect 932 -274 966 -240
rect 1128 -274 1162 -240
rect 1324 -274 1358 -240
rect 1520 -274 1554 -240
rect 1716 -274 1750 -240
rect 1912 -274 1946 -240
rect 2108 -274 2142 -240
rect 2304 -274 2338 -240
rect 2500 -274 2534 -240
rect 2696 -274 2730 -240
rect 2892 -274 2926 -240
rect 638 -784 672 -750
rect 834 -784 868 -750
rect 1030 -784 1064 -750
rect 1226 -784 1260 -750
rect 1422 -784 1456 -750
rect 1618 -784 1652 -750
rect 1814 -784 1848 -750
rect 2010 -784 2044 -750
rect 2206 -784 2240 -750
rect 2402 -784 2436 -750
rect 2598 -784 2632 -750
rect 2794 -784 2828 -750
rect 2990 -784 3024 -750
rect 639 -892 673 -858
rect 835 -892 869 -858
rect 1031 -892 1065 -858
rect 1227 -892 1261 -858
rect 1423 -892 1457 -858
rect 1619 -892 1653 -858
rect 1815 -892 1849 -858
rect 2011 -892 2045 -858
rect 2207 -892 2241 -858
rect 2403 -892 2437 -858
rect 2599 -892 2633 -858
rect 2795 -892 2829 -858
rect 2991 -892 3025 -858
rect 737 -1402 771 -1368
rect 933 -1402 967 -1368
rect 1129 -1402 1163 -1368
rect 1325 -1402 1359 -1368
rect 1521 -1402 1555 -1368
rect 1717 -1402 1751 -1368
rect 1913 -1402 1947 -1368
rect 2109 -1402 2143 -1368
rect 2305 -1402 2339 -1368
rect 2501 -1402 2535 -1368
rect 2697 -1402 2731 -1368
rect 2893 -1402 2927 -1368
rect 736 -1718 770 -1684
rect 932 -1718 966 -1684
rect 1128 -1718 1162 -1684
rect 1324 -1718 1358 -1684
rect 1520 -1718 1554 -1684
rect 1716 -1718 1750 -1684
rect 1912 -1718 1946 -1684
rect 2108 -1718 2142 -1684
rect 2304 -1718 2338 -1684
rect 2500 -1718 2534 -1684
rect 2696 -1718 2730 -1684
rect 2892 -1718 2926 -1684
rect 638 -2228 672 -2194
rect 834 -2228 868 -2194
rect 1030 -2228 1064 -2194
rect 1226 -2228 1260 -2194
rect 1422 -2228 1456 -2194
rect 1618 -2228 1652 -2194
rect 1814 -2228 1848 -2194
rect 2010 -2228 2044 -2194
rect 2206 -2228 2240 -2194
rect 2402 -2228 2436 -2194
rect 2598 -2228 2632 -2194
rect 2794 -2228 2828 -2194
rect 2990 -2228 3024 -2194
rect 639 -2336 673 -2302
rect 835 -2336 869 -2302
rect 1031 -2336 1065 -2302
rect 1227 -2336 1261 -2302
rect 1423 -2336 1457 -2302
rect 1619 -2336 1653 -2302
rect 1815 -2336 1849 -2302
rect 2011 -2336 2045 -2302
rect 2207 -2336 2241 -2302
rect 2403 -2336 2437 -2302
rect 2599 -2336 2633 -2302
rect 2795 -2336 2829 -2302
rect 2991 -2336 3025 -2302
rect 737 -2846 771 -2812
rect 933 -2846 967 -2812
rect 1129 -2846 1163 -2812
rect 1325 -2846 1359 -2812
rect 1521 -2846 1555 -2812
rect 1717 -2846 1751 -2812
rect 1913 -2846 1947 -2812
rect 2109 -2846 2143 -2812
rect 2305 -2846 2339 -2812
rect 2501 -2846 2535 -2812
rect 2697 -2846 2731 -2812
rect 2893 -2846 2927 -2812
<< metal1 >>
rect 623 1236 2061 1252
rect 623 1202 737 1236
rect 771 1202 933 1236
rect 967 1202 1129 1236
rect 1163 1202 1325 1236
rect 1359 1202 1521 1236
rect 1555 1202 1717 1236
rect 1751 1202 1913 1236
rect 1947 1202 2061 1236
rect 623 1186 2061 1202
rect 2421 1236 3859 1252
rect 2421 1202 2535 1236
rect 2569 1202 2731 1236
rect 2765 1202 2927 1236
rect 2961 1202 3123 1236
rect 3157 1202 3319 1236
rect 3353 1202 3515 1236
rect 3549 1202 3711 1236
rect 3745 1202 3859 1236
rect 2421 1186 3859 1202
rect 669 995 679 1155
rect 731 995 741 1155
rect 865 995 875 1155
rect 927 995 937 1155
rect 1061 995 1071 1155
rect 1123 995 1133 1155
rect 1257 995 1267 1155
rect 1319 995 1329 1155
rect 1453 995 1463 1155
rect 1515 995 1525 1155
rect 1649 995 1659 1155
rect 1711 995 1721 1155
rect 1845 995 1855 1155
rect 1907 995 1917 1155
rect 2041 995 2051 1155
rect 2103 995 2113 1155
rect 2467 995 2477 1155
rect 2529 995 2539 1155
rect 2663 995 2673 1155
rect 2725 995 2735 1155
rect 2859 995 2869 1155
rect 2921 995 2931 1155
rect 3055 995 3065 1155
rect 3117 995 3127 1155
rect 3251 995 3261 1155
rect 3313 995 3323 1155
rect 3447 995 3457 1155
rect 3509 995 3519 1155
rect 3643 995 3653 1155
rect 3705 995 3715 1155
rect 3839 995 3849 1155
rect 3901 995 3911 1155
rect 571 755 581 915
rect 633 755 643 915
rect 767 755 777 915
rect 829 755 839 915
rect 963 755 973 915
rect 1025 755 1035 915
rect 1159 755 1169 915
rect 1221 755 1231 915
rect 1355 755 1365 915
rect 1417 755 1427 915
rect 1551 755 1561 915
rect 1613 755 1623 915
rect 1747 755 1757 915
rect 1809 755 1819 915
rect 1943 755 1953 915
rect 2005 755 2015 915
rect 2369 755 2379 915
rect 2431 755 2441 915
rect 2565 755 2575 915
rect 2627 755 2637 915
rect 2761 755 2771 915
rect 2823 755 2833 915
rect 2957 755 2967 915
rect 3019 755 3029 915
rect 3153 755 3163 915
rect 3215 755 3225 915
rect 3349 755 3359 915
rect 3411 755 3421 915
rect 3545 755 3555 915
rect 3607 755 3617 915
rect 3741 755 3751 915
rect 3803 755 3813 915
rect 623 708 2061 724
rect 623 674 639 708
rect 673 674 835 708
rect 869 674 1031 708
rect 1065 674 1227 708
rect 1261 674 1423 708
rect 1457 674 1619 708
rect 1653 674 1815 708
rect 1849 674 2011 708
rect 2045 674 2061 708
rect 623 658 2061 674
rect 2421 708 3859 724
rect 2421 674 2437 708
rect 2471 674 2633 708
rect 2667 674 2829 708
rect 2863 674 3025 708
rect 3059 674 3221 708
rect 3255 674 3417 708
rect 3451 674 3613 708
rect 3647 674 3809 708
rect 3843 674 3859 708
rect 2421 658 3859 674
rect 623 600 2061 616
rect 623 566 639 600
rect 673 566 835 600
rect 869 566 1031 600
rect 1065 566 1227 600
rect 1261 566 1423 600
rect 1457 566 1619 600
rect 1653 566 1815 600
rect 1849 566 2011 600
rect 2045 566 2061 600
rect 623 550 2061 566
rect 2421 600 3859 616
rect 2421 566 2437 600
rect 2471 566 2633 600
rect 2667 566 2829 600
rect 2863 566 3025 600
rect 3059 566 3221 600
rect 3255 566 3417 600
rect 3451 566 3613 600
rect 3647 566 3809 600
rect 3843 566 3859 600
rect 2421 550 3859 566
rect 571 359 581 519
rect 633 359 643 519
rect 767 359 777 519
rect 829 359 839 519
rect 963 359 973 519
rect 1025 359 1035 519
rect 1159 359 1169 519
rect 1221 359 1231 519
rect 1355 359 1365 519
rect 1417 359 1427 519
rect 1551 359 1561 519
rect 1613 359 1623 519
rect 1747 359 1757 519
rect 1809 359 1819 519
rect 1943 359 1953 519
rect 2005 359 2015 519
rect 2369 359 2379 519
rect 2431 359 2441 519
rect 2565 359 2575 519
rect 2627 359 2637 519
rect 2761 359 2771 519
rect 2823 359 2833 519
rect 2957 359 2967 519
rect 3019 359 3029 519
rect 3153 359 3163 519
rect 3215 359 3225 519
rect 3349 359 3359 519
rect 3411 359 3421 519
rect 3545 359 3555 519
rect 3607 359 3617 519
rect 3741 359 3751 519
rect 3803 359 3813 519
rect 669 119 679 279
rect 731 119 741 279
rect 865 119 875 279
rect 927 119 937 279
rect 1061 119 1071 279
rect 1123 119 1133 279
rect 1257 119 1267 279
rect 1319 119 1329 279
rect 1453 119 1463 279
rect 1515 119 1525 279
rect 1649 119 1659 279
rect 1711 119 1721 279
rect 1845 119 1855 279
rect 1907 119 1917 279
rect 2041 119 2051 279
rect 2103 119 2113 279
rect 2467 119 2477 279
rect 2529 119 2539 279
rect 2663 119 2673 279
rect 2725 119 2735 279
rect 2859 119 2869 279
rect 2921 119 2931 279
rect 3055 119 3065 279
rect 3117 119 3127 279
rect 3251 119 3261 279
rect 3313 119 3323 279
rect 3447 119 3457 279
rect 3509 119 3519 279
rect 3643 119 3653 279
rect 3705 119 3715 279
rect 3839 119 3849 279
rect 3901 119 3911 279
rect 623 72 2061 88
rect 623 38 737 72
rect 771 38 933 72
rect 967 38 1129 72
rect 1163 38 1325 72
rect 1359 38 1521 72
rect 1555 38 1717 72
rect 1751 38 1913 72
rect 1947 38 2061 72
rect 623 22 2061 38
rect 2421 72 3859 88
rect 2421 38 2535 72
rect 2569 38 2731 72
rect 2765 38 2927 72
rect 2961 38 3123 72
rect 3157 38 3319 72
rect 3353 38 3515 72
rect 3549 38 3711 72
rect 3745 38 3859 72
rect 2421 22 3859 38
rect 622 -240 3040 -224
rect 622 -274 736 -240
rect 770 -274 932 -240
rect 966 -274 1128 -240
rect 1162 -274 1324 -240
rect 1358 -274 1520 -240
rect 1554 -274 1716 -240
rect 1750 -274 1912 -240
rect 1946 -274 2108 -240
rect 2142 -274 2304 -240
rect 2338 -274 2500 -240
rect 2534 -274 2696 -240
rect 2730 -274 2892 -240
rect 2926 -274 3040 -240
rect 622 -284 3040 -274
rect 669 -472 679 -312
rect 731 -472 741 -312
rect 865 -472 875 -312
rect 927 -472 937 -312
rect 1061 -472 1071 -312
rect 1123 -472 1133 -312
rect 1257 -472 1267 -312
rect 1319 -472 1329 -312
rect 1453 -472 1463 -312
rect 1515 -472 1525 -312
rect 1649 -472 1659 -312
rect 1711 -472 1721 -312
rect 1845 -472 1855 -312
rect 1907 -472 1917 -312
rect 2041 -472 2051 -312
rect 2103 -472 2113 -312
rect 2237 -472 2247 -312
rect 2299 -472 2309 -312
rect 2433 -472 2443 -312
rect 2495 -472 2505 -312
rect 2629 -472 2639 -312
rect 2691 -472 2701 -312
rect 2825 -472 2835 -312
rect 2887 -472 2897 -312
rect 3021 -472 3031 -312
rect 3083 -472 3093 -312
rect 571 -712 581 -552
rect 633 -712 643 -552
rect 767 -712 777 -552
rect 829 -712 839 -552
rect 963 -712 973 -552
rect 1025 -712 1035 -552
rect 1159 -712 1169 -552
rect 1221 -712 1231 -552
rect 1355 -712 1365 -552
rect 1417 -712 1427 -552
rect 1551 -712 1561 -552
rect 1613 -712 1623 -552
rect 1747 -712 1757 -552
rect 1809 -712 1819 -552
rect 1943 -712 1953 -552
rect 2005 -712 2015 -552
rect 2139 -712 2149 -552
rect 2201 -712 2211 -552
rect 2335 -712 2345 -552
rect 2397 -712 2407 -552
rect 2531 -712 2541 -552
rect 2593 -712 2603 -552
rect 2727 -712 2737 -552
rect 2789 -712 2799 -552
rect 2923 -712 2933 -552
rect 2985 -712 2995 -552
rect 622 -750 3040 -740
rect 622 -784 638 -750
rect 672 -784 834 -750
rect 868 -784 1030 -750
rect 1064 -784 1226 -750
rect 1260 -784 1422 -750
rect 1456 -784 1618 -750
rect 1652 -784 1814 -750
rect 1848 -784 2010 -750
rect 2044 -784 2206 -750
rect 2240 -784 2402 -750
rect 2436 -784 2598 -750
rect 2632 -784 2794 -750
rect 2828 -784 2990 -750
rect 3024 -784 3040 -750
rect 622 -800 3040 -784
rect 623 -858 3041 -842
rect 623 -892 639 -858
rect 673 -892 835 -858
rect 869 -892 1031 -858
rect 1065 -892 1227 -858
rect 1261 -892 1423 -858
rect 1457 -892 1619 -858
rect 1653 -892 1815 -858
rect 1849 -892 2011 -858
rect 2045 -892 2207 -858
rect 2241 -892 2403 -858
rect 2437 -892 2599 -858
rect 2633 -892 2795 -858
rect 2829 -892 2991 -858
rect 3025 -892 3041 -858
rect 623 -902 3041 -892
rect 571 -1090 581 -930
rect 633 -1090 643 -930
rect 767 -1090 777 -930
rect 829 -1090 839 -930
rect 963 -1090 973 -930
rect 1025 -1090 1035 -930
rect 1159 -1090 1169 -930
rect 1221 -1090 1231 -930
rect 1355 -1090 1365 -930
rect 1417 -1090 1427 -930
rect 1551 -1090 1561 -930
rect 1613 -1090 1623 -930
rect 1747 -1090 1757 -930
rect 1809 -1090 1819 -930
rect 1943 -1090 1953 -930
rect 2005 -1090 2015 -930
rect 2139 -1090 2149 -930
rect 2201 -1090 2211 -930
rect 2335 -1090 2345 -930
rect 2397 -1090 2407 -930
rect 2531 -1090 2541 -930
rect 2593 -1090 2603 -930
rect 2727 -1090 2737 -930
rect 2789 -1090 2799 -930
rect 2923 -1090 2933 -930
rect 2985 -1090 2995 -930
rect 669 -1330 679 -1170
rect 731 -1330 741 -1170
rect 865 -1330 875 -1170
rect 927 -1330 937 -1170
rect 1061 -1330 1071 -1170
rect 1123 -1330 1133 -1170
rect 1257 -1330 1267 -1170
rect 1319 -1330 1329 -1170
rect 1453 -1330 1463 -1170
rect 1515 -1330 1525 -1170
rect 1649 -1330 1659 -1170
rect 1711 -1330 1721 -1170
rect 1845 -1330 1855 -1170
rect 1907 -1330 1917 -1170
rect 2041 -1330 2051 -1170
rect 2103 -1330 2113 -1170
rect 2237 -1330 2247 -1170
rect 2299 -1330 2309 -1170
rect 2433 -1330 2443 -1170
rect 2495 -1330 2505 -1170
rect 2629 -1330 2639 -1170
rect 2691 -1330 2701 -1170
rect 2825 -1330 2835 -1170
rect 2887 -1330 2897 -1170
rect 3021 -1330 3031 -1170
rect 3083 -1330 3093 -1170
rect 623 -1368 3041 -1358
rect 623 -1402 737 -1368
rect 771 -1402 933 -1368
rect 967 -1402 1129 -1368
rect 1163 -1402 1325 -1368
rect 1359 -1402 1521 -1368
rect 1555 -1402 1717 -1368
rect 1751 -1402 1913 -1368
rect 1947 -1402 2109 -1368
rect 2143 -1402 2305 -1368
rect 2339 -1402 2501 -1368
rect 2535 -1402 2697 -1368
rect 2731 -1402 2893 -1368
rect 2927 -1402 3041 -1368
rect 623 -1418 3041 -1402
rect 622 -1684 3040 -1668
rect 622 -1718 736 -1684
rect 770 -1718 932 -1684
rect 966 -1718 1128 -1684
rect 1162 -1718 1324 -1684
rect 1358 -1718 1520 -1684
rect 1554 -1718 1716 -1684
rect 1750 -1718 1912 -1684
rect 1946 -1718 2108 -1684
rect 2142 -1718 2304 -1684
rect 2338 -1718 2500 -1684
rect 2534 -1718 2696 -1684
rect 2730 -1718 2892 -1684
rect 2926 -1718 3040 -1684
rect 622 -1728 3040 -1718
rect 669 -1916 679 -1756
rect 731 -1916 741 -1756
rect 865 -1916 875 -1756
rect 927 -1916 937 -1756
rect 1061 -1916 1071 -1756
rect 1123 -1916 1133 -1756
rect 1257 -1916 1267 -1756
rect 1319 -1916 1329 -1756
rect 1453 -1916 1463 -1756
rect 1515 -1916 1525 -1756
rect 1649 -1916 1659 -1756
rect 1711 -1916 1721 -1756
rect 1845 -1916 1855 -1756
rect 1907 -1916 1917 -1756
rect 2041 -1916 2051 -1756
rect 2103 -1916 2113 -1756
rect 2237 -1916 2247 -1756
rect 2299 -1916 2309 -1756
rect 2433 -1916 2443 -1756
rect 2495 -1916 2505 -1756
rect 2629 -1916 2639 -1756
rect 2691 -1916 2701 -1756
rect 2825 -1916 2835 -1756
rect 2887 -1916 2897 -1756
rect 3021 -1916 3031 -1756
rect 3083 -1916 3093 -1756
rect 571 -2156 581 -1996
rect 633 -2156 643 -1996
rect 767 -2156 777 -1996
rect 829 -2156 839 -1996
rect 963 -2156 973 -1996
rect 1025 -2156 1035 -1996
rect 1159 -2156 1169 -1996
rect 1221 -2156 1231 -1996
rect 1355 -2156 1365 -1996
rect 1417 -2156 1427 -1996
rect 1551 -2156 1561 -1996
rect 1613 -2156 1623 -1996
rect 1747 -2156 1757 -1996
rect 1809 -2156 1819 -1996
rect 1943 -2156 1953 -1996
rect 2005 -2156 2015 -1996
rect 2139 -2156 2149 -1996
rect 2201 -2156 2211 -1996
rect 2335 -2156 2345 -1996
rect 2397 -2156 2407 -1996
rect 2531 -2156 2541 -1996
rect 2593 -2156 2603 -1996
rect 2727 -2156 2737 -1996
rect 2789 -2156 2799 -1996
rect 2923 -2156 2933 -1996
rect 2985 -2156 2995 -1996
rect 622 -2194 3040 -2184
rect 622 -2228 638 -2194
rect 672 -2228 834 -2194
rect 868 -2228 1030 -2194
rect 1064 -2228 1226 -2194
rect 1260 -2228 1422 -2194
rect 1456 -2228 1618 -2194
rect 1652 -2228 1814 -2194
rect 1848 -2228 2010 -2194
rect 2044 -2228 2206 -2194
rect 2240 -2228 2402 -2194
rect 2436 -2228 2598 -2194
rect 2632 -2228 2794 -2194
rect 2828 -2228 2990 -2194
rect 3024 -2228 3040 -2194
rect 622 -2244 3040 -2228
rect 623 -2302 3041 -2286
rect 623 -2336 639 -2302
rect 673 -2336 835 -2302
rect 869 -2336 1031 -2302
rect 1065 -2336 1227 -2302
rect 1261 -2336 1423 -2302
rect 1457 -2336 1619 -2302
rect 1653 -2336 1815 -2302
rect 1849 -2336 2011 -2302
rect 2045 -2336 2207 -2302
rect 2241 -2336 2403 -2302
rect 2437 -2336 2599 -2302
rect 2633 -2336 2795 -2302
rect 2829 -2336 2991 -2302
rect 3025 -2336 3041 -2302
rect 623 -2346 3041 -2336
rect 571 -2534 581 -2374
rect 633 -2534 643 -2374
rect 767 -2534 777 -2374
rect 829 -2534 839 -2374
rect 963 -2534 973 -2374
rect 1025 -2534 1035 -2374
rect 1159 -2534 1169 -2374
rect 1221 -2534 1231 -2374
rect 1355 -2534 1365 -2374
rect 1417 -2534 1427 -2374
rect 1551 -2534 1561 -2374
rect 1613 -2534 1623 -2374
rect 1747 -2534 1757 -2374
rect 1809 -2534 1819 -2374
rect 1943 -2534 1953 -2374
rect 2005 -2534 2015 -2374
rect 2139 -2534 2149 -2374
rect 2201 -2534 2211 -2374
rect 2335 -2534 2345 -2374
rect 2397 -2534 2407 -2374
rect 2531 -2534 2541 -2374
rect 2593 -2534 2603 -2374
rect 2727 -2534 2737 -2374
rect 2789 -2534 2799 -2374
rect 2923 -2534 2933 -2374
rect 2985 -2534 2995 -2374
rect 669 -2774 679 -2614
rect 731 -2774 741 -2614
rect 865 -2774 875 -2614
rect 927 -2774 937 -2614
rect 1061 -2774 1071 -2614
rect 1123 -2774 1133 -2614
rect 1257 -2774 1267 -2614
rect 1319 -2774 1329 -2614
rect 1453 -2774 1463 -2614
rect 1515 -2774 1525 -2614
rect 1649 -2774 1659 -2614
rect 1711 -2774 1721 -2614
rect 1845 -2774 1855 -2614
rect 1907 -2774 1917 -2614
rect 2041 -2774 2051 -2614
rect 2103 -2774 2113 -2614
rect 2237 -2774 2247 -2614
rect 2299 -2774 2309 -2614
rect 2433 -2774 2443 -2614
rect 2495 -2774 2505 -2614
rect 2629 -2774 2639 -2614
rect 2691 -2774 2701 -2614
rect 2825 -2774 2835 -2614
rect 2887 -2774 2897 -2614
rect 3021 -2774 3031 -2614
rect 3083 -2774 3093 -2614
rect 623 -2812 3041 -2802
rect 623 -2846 737 -2812
rect 771 -2846 933 -2812
rect 967 -2846 1129 -2812
rect 1163 -2846 1325 -2812
rect 1359 -2846 1521 -2812
rect 1555 -2846 1717 -2812
rect 1751 -2846 1913 -2812
rect 1947 -2846 2109 -2812
rect 2143 -2846 2305 -2812
rect 2339 -2846 2501 -2812
rect 2535 -2846 2697 -2812
rect 2731 -2846 2893 -2812
rect 2927 -2846 3041 -2812
rect 623 -2862 3041 -2846
<< via1 >>
rect 679 995 731 1155
rect 875 995 927 1155
rect 1071 995 1123 1155
rect 1267 995 1319 1155
rect 1463 995 1515 1155
rect 1659 995 1711 1155
rect 1855 995 1907 1155
rect 2051 995 2103 1155
rect 2477 995 2529 1155
rect 2673 995 2725 1155
rect 2869 995 2921 1155
rect 3065 995 3117 1155
rect 3261 995 3313 1155
rect 3457 995 3509 1155
rect 3653 995 3705 1155
rect 3849 995 3901 1155
rect 581 755 633 915
rect 777 755 829 915
rect 973 755 1025 915
rect 1169 755 1221 915
rect 1365 755 1417 915
rect 1561 755 1613 915
rect 1757 755 1809 915
rect 1953 755 2005 915
rect 2379 755 2431 915
rect 2575 755 2627 915
rect 2771 755 2823 915
rect 2967 755 3019 915
rect 3163 755 3215 915
rect 3359 755 3411 915
rect 3555 755 3607 915
rect 3751 755 3803 915
rect 581 359 633 519
rect 777 359 829 519
rect 973 359 1025 519
rect 1169 359 1221 519
rect 1365 359 1417 519
rect 1561 359 1613 519
rect 1757 359 1809 519
rect 1953 359 2005 519
rect 2379 359 2431 519
rect 2575 359 2627 519
rect 2771 359 2823 519
rect 2967 359 3019 519
rect 3163 359 3215 519
rect 3359 359 3411 519
rect 3555 359 3607 519
rect 3751 359 3803 519
rect 679 119 731 279
rect 875 119 927 279
rect 1071 119 1123 279
rect 1267 119 1319 279
rect 1463 119 1515 279
rect 1659 119 1711 279
rect 1855 119 1907 279
rect 2051 119 2103 279
rect 2477 119 2529 279
rect 2673 119 2725 279
rect 2869 119 2921 279
rect 3065 119 3117 279
rect 3261 119 3313 279
rect 3457 119 3509 279
rect 3653 119 3705 279
rect 3849 119 3901 279
rect 679 -472 731 -312
rect 875 -472 927 -312
rect 1071 -472 1123 -312
rect 1267 -472 1319 -312
rect 1463 -472 1515 -312
rect 1659 -472 1711 -312
rect 1855 -472 1907 -312
rect 2051 -472 2103 -312
rect 2247 -472 2299 -312
rect 2443 -472 2495 -312
rect 2639 -472 2691 -312
rect 2835 -472 2887 -312
rect 3031 -472 3083 -312
rect 581 -712 633 -552
rect 777 -712 829 -552
rect 973 -712 1025 -552
rect 1169 -712 1221 -552
rect 1365 -712 1417 -552
rect 1561 -712 1613 -552
rect 1757 -712 1809 -552
rect 1953 -712 2005 -552
rect 2149 -712 2201 -552
rect 2345 -712 2397 -552
rect 2541 -712 2593 -552
rect 2737 -712 2789 -552
rect 2933 -712 2985 -552
rect 581 -1090 633 -930
rect 777 -1090 829 -930
rect 973 -1090 1025 -930
rect 1169 -1090 1221 -930
rect 1365 -1090 1417 -930
rect 1561 -1090 1613 -930
rect 1757 -1090 1809 -930
rect 1953 -1090 2005 -930
rect 2149 -1090 2201 -930
rect 2345 -1090 2397 -930
rect 2541 -1090 2593 -930
rect 2737 -1090 2789 -930
rect 2933 -1090 2985 -930
rect 679 -1330 731 -1170
rect 875 -1330 927 -1170
rect 1071 -1330 1123 -1170
rect 1267 -1330 1319 -1170
rect 1463 -1330 1515 -1170
rect 1659 -1330 1711 -1170
rect 1855 -1330 1907 -1170
rect 2051 -1330 2103 -1170
rect 2247 -1330 2299 -1170
rect 2443 -1330 2495 -1170
rect 2639 -1330 2691 -1170
rect 2835 -1330 2887 -1170
rect 3031 -1330 3083 -1170
rect 679 -1916 731 -1756
rect 875 -1916 927 -1756
rect 1071 -1916 1123 -1756
rect 1267 -1916 1319 -1756
rect 1463 -1916 1515 -1756
rect 1659 -1916 1711 -1756
rect 1855 -1916 1907 -1756
rect 2051 -1916 2103 -1756
rect 2247 -1916 2299 -1756
rect 2443 -1916 2495 -1756
rect 2639 -1916 2691 -1756
rect 2835 -1916 2887 -1756
rect 3031 -1916 3083 -1756
rect 581 -2156 633 -1996
rect 777 -2156 829 -1996
rect 973 -2156 1025 -1996
rect 1169 -2156 1221 -1996
rect 1365 -2156 1417 -1996
rect 1561 -2156 1613 -1996
rect 1757 -2156 1809 -1996
rect 1953 -2156 2005 -1996
rect 2149 -2156 2201 -1996
rect 2345 -2156 2397 -1996
rect 2541 -2156 2593 -1996
rect 2737 -2156 2789 -1996
rect 2933 -2156 2985 -1996
rect 581 -2534 633 -2374
rect 777 -2534 829 -2374
rect 973 -2534 1025 -2374
rect 1169 -2534 1221 -2374
rect 1365 -2534 1417 -2374
rect 1561 -2534 1613 -2374
rect 1757 -2534 1809 -2374
rect 1953 -2534 2005 -2374
rect 2149 -2534 2201 -2374
rect 2345 -2534 2397 -2374
rect 2541 -2534 2593 -2374
rect 2737 -2534 2789 -2374
rect 2933 -2534 2985 -2374
rect 679 -2774 731 -2614
rect 875 -2774 927 -2614
rect 1071 -2774 1123 -2614
rect 1267 -2774 1319 -2614
rect 1463 -2774 1515 -2614
rect 1659 -2774 1711 -2614
rect 1855 -2774 1907 -2614
rect 2051 -2774 2103 -2614
rect 2247 -2774 2299 -2614
rect 2443 -2774 2495 -2614
rect 2639 -2774 2691 -2614
rect 2835 -2774 2887 -2614
rect 3031 -2774 3083 -2614
<< metal2 >>
rect 679 1155 731 1165
rect 679 985 731 995
rect 875 1155 927 1165
rect 875 985 927 995
rect 1071 1155 1123 1165
rect 1071 985 1123 995
rect 1267 1155 1319 1165
rect 1267 985 1319 995
rect 1463 1155 1515 1165
rect 1463 985 1515 995
rect 1659 1155 1711 1165
rect 1659 985 1711 995
rect 1855 1155 1907 1165
rect 1855 985 1907 995
rect 2051 1155 2103 1165
rect 2051 985 2103 995
rect 2477 1155 2529 1165
rect 2477 985 2529 995
rect 2673 1155 2725 1165
rect 2673 985 2725 995
rect 2869 1155 2921 1165
rect 2869 985 2921 995
rect 3065 1155 3117 1165
rect 3065 985 3117 995
rect 3261 1155 3313 1165
rect 3261 985 3313 995
rect 3457 1155 3509 1165
rect 3457 985 3509 995
rect 3653 1155 3705 1165
rect 3653 985 3705 995
rect 3849 1155 3901 1165
rect 3849 985 3901 995
rect 581 915 633 925
rect 581 745 633 755
rect 777 915 829 925
rect 777 745 829 755
rect 973 915 1025 925
rect 973 745 1025 755
rect 1169 915 1221 925
rect 1169 745 1221 755
rect 1365 915 1417 925
rect 1365 745 1417 755
rect 1561 915 1613 925
rect 1561 745 1613 755
rect 1757 915 1809 925
rect 1757 745 1809 755
rect 1953 915 2005 925
rect 1953 745 2005 755
rect 2379 915 2431 925
rect 2379 745 2431 755
rect 2575 915 2627 925
rect 2575 745 2627 755
rect 2771 915 2823 925
rect 2771 745 2823 755
rect 2967 915 3019 925
rect 2967 745 3019 755
rect 3163 915 3215 925
rect 3163 745 3215 755
rect 3359 915 3411 925
rect 3359 745 3411 755
rect 3555 915 3607 925
rect 3555 745 3607 755
rect 3751 915 3803 925
rect 3751 745 3803 755
rect 581 519 633 529
rect 581 349 633 359
rect 777 519 829 529
rect 777 349 829 359
rect 973 519 1025 529
rect 973 349 1025 359
rect 1169 519 1221 529
rect 1169 349 1221 359
rect 1365 519 1417 529
rect 1365 349 1417 359
rect 1561 519 1613 529
rect 1561 349 1613 359
rect 1757 519 1809 529
rect 1757 349 1809 359
rect 1953 519 2005 529
rect 1953 349 2005 359
rect 2379 519 2431 529
rect 2379 349 2431 359
rect 2575 519 2627 529
rect 2575 349 2627 359
rect 2771 519 2823 529
rect 2771 349 2823 359
rect 2967 519 3019 529
rect 2967 349 3019 359
rect 3163 519 3215 529
rect 3163 349 3215 359
rect 3359 519 3411 529
rect 3359 349 3411 359
rect 3555 519 3607 529
rect 3555 349 3607 359
rect 3751 519 3803 529
rect 3751 349 3803 359
rect 679 279 731 289
rect 679 109 731 119
rect 875 279 927 289
rect 875 109 927 119
rect 1071 279 1123 289
rect 1071 109 1123 119
rect 1267 279 1319 289
rect 1267 109 1319 119
rect 1463 279 1515 289
rect 1463 109 1515 119
rect 1659 279 1711 289
rect 1659 109 1711 119
rect 1855 279 1907 289
rect 1855 109 1907 119
rect 2051 279 2103 289
rect 2051 109 2103 119
rect 2477 279 2529 289
rect 2477 109 2529 119
rect 2673 279 2725 289
rect 2673 109 2725 119
rect 2869 279 2921 289
rect 2869 109 2921 119
rect 3065 279 3117 289
rect 3065 109 3117 119
rect 3261 279 3313 289
rect 3261 109 3313 119
rect 3457 279 3509 289
rect 3457 109 3509 119
rect 3653 279 3705 289
rect 3653 109 3705 119
rect 3849 279 3901 289
rect 3849 109 3901 119
rect 679 -312 731 -302
rect 679 -482 731 -472
rect 875 -312 927 -302
rect 875 -482 927 -472
rect 1071 -312 1123 -302
rect 1071 -482 1123 -472
rect 1267 -312 1319 -302
rect 1267 -482 1319 -472
rect 1463 -312 1515 -302
rect 1463 -482 1515 -472
rect 1659 -312 1711 -302
rect 1659 -482 1711 -472
rect 1855 -312 1907 -302
rect 1855 -482 1907 -472
rect 2051 -312 2103 -302
rect 2051 -482 2103 -472
rect 2247 -312 2299 -302
rect 2247 -482 2299 -472
rect 2443 -312 2495 -302
rect 2443 -482 2495 -472
rect 2639 -312 2691 -302
rect 2639 -482 2691 -472
rect 2835 -312 2887 -302
rect 2835 -482 2887 -472
rect 3031 -312 3083 -302
rect 3031 -482 3083 -472
rect 581 -552 633 -542
rect 581 -722 633 -712
rect 777 -552 829 -542
rect 777 -722 829 -712
rect 973 -552 1025 -542
rect 973 -722 1025 -712
rect 1169 -552 1221 -542
rect 1169 -722 1221 -712
rect 1365 -552 1417 -542
rect 1365 -722 1417 -712
rect 1561 -552 1613 -542
rect 1561 -722 1613 -712
rect 1757 -552 1809 -542
rect 1757 -722 1809 -712
rect 1953 -552 2005 -542
rect 1953 -722 2005 -712
rect 2149 -552 2201 -542
rect 2149 -722 2201 -712
rect 2345 -552 2397 -542
rect 2345 -722 2397 -712
rect 2541 -552 2593 -542
rect 2541 -722 2593 -712
rect 2737 -552 2789 -542
rect 2737 -722 2789 -712
rect 2933 -552 2985 -542
rect 2933 -722 2985 -712
rect 581 -930 633 -920
rect 581 -1100 633 -1090
rect 777 -930 829 -920
rect 777 -1100 829 -1090
rect 973 -930 1025 -920
rect 973 -1100 1025 -1090
rect 1169 -930 1221 -920
rect 1169 -1100 1221 -1090
rect 1365 -930 1417 -920
rect 1365 -1100 1417 -1090
rect 1561 -930 1613 -920
rect 1561 -1100 1613 -1090
rect 1757 -930 1809 -920
rect 1757 -1100 1809 -1090
rect 1953 -930 2005 -920
rect 1953 -1100 2005 -1090
rect 2149 -930 2201 -920
rect 2149 -1100 2201 -1090
rect 2345 -930 2397 -920
rect 2345 -1100 2397 -1090
rect 2541 -930 2593 -920
rect 2541 -1100 2593 -1090
rect 2737 -930 2789 -920
rect 2737 -1100 2789 -1090
rect 2933 -930 2985 -920
rect 2933 -1100 2985 -1090
rect 679 -1170 731 -1160
rect 679 -1340 731 -1330
rect 875 -1170 927 -1160
rect 875 -1340 927 -1330
rect 1071 -1170 1123 -1160
rect 1071 -1340 1123 -1330
rect 1267 -1170 1319 -1160
rect 1267 -1340 1319 -1330
rect 1463 -1170 1515 -1160
rect 1463 -1340 1515 -1330
rect 1659 -1170 1711 -1160
rect 1659 -1340 1711 -1330
rect 1855 -1170 1907 -1160
rect 1855 -1340 1907 -1330
rect 2051 -1170 2103 -1160
rect 2051 -1340 2103 -1330
rect 2247 -1170 2299 -1160
rect 2247 -1340 2299 -1330
rect 2443 -1170 2495 -1160
rect 2443 -1340 2495 -1330
rect 2639 -1170 2691 -1160
rect 2639 -1340 2691 -1330
rect 2835 -1170 2887 -1160
rect 2835 -1340 2887 -1330
rect 3031 -1170 3083 -1160
rect 3031 -1340 3083 -1330
rect 679 -1756 731 -1746
rect 679 -1926 731 -1916
rect 875 -1756 927 -1746
rect 875 -1926 927 -1916
rect 1071 -1756 1123 -1746
rect 1071 -1926 1123 -1916
rect 1267 -1756 1319 -1746
rect 1267 -1926 1319 -1916
rect 1463 -1756 1515 -1746
rect 1463 -1926 1515 -1916
rect 1659 -1756 1711 -1746
rect 1659 -1926 1711 -1916
rect 1855 -1756 1907 -1746
rect 1855 -1926 1907 -1916
rect 2051 -1756 2103 -1746
rect 2051 -1926 2103 -1916
rect 2247 -1756 2299 -1746
rect 2247 -1926 2299 -1916
rect 2443 -1756 2495 -1746
rect 2443 -1926 2495 -1916
rect 2639 -1756 2691 -1746
rect 2639 -1926 2691 -1916
rect 2835 -1756 2887 -1746
rect 2835 -1926 2887 -1916
rect 3031 -1756 3083 -1746
rect 3031 -1926 3083 -1916
rect 581 -1996 633 -1986
rect 581 -2166 633 -2156
rect 777 -1996 829 -1986
rect 777 -2166 829 -2156
rect 973 -1996 1025 -1986
rect 973 -2166 1025 -2156
rect 1169 -1996 1221 -1986
rect 1169 -2166 1221 -2156
rect 1365 -1996 1417 -1986
rect 1365 -2166 1417 -2156
rect 1561 -1996 1613 -1986
rect 1561 -2166 1613 -2156
rect 1757 -1996 1809 -1986
rect 1757 -2166 1809 -2156
rect 1953 -1996 2005 -1986
rect 1953 -2166 2005 -2156
rect 2149 -1996 2201 -1986
rect 2149 -2166 2201 -2156
rect 2345 -1996 2397 -1986
rect 2345 -2166 2397 -2156
rect 2541 -1996 2593 -1986
rect 2541 -2166 2593 -2156
rect 2737 -1996 2789 -1986
rect 2737 -2166 2789 -2156
rect 2933 -1996 2985 -1986
rect 2933 -2166 2985 -2156
rect 581 -2374 633 -2364
rect 581 -2544 633 -2534
rect 777 -2374 829 -2364
rect 777 -2544 829 -2534
rect 973 -2374 1025 -2364
rect 973 -2544 1025 -2534
rect 1169 -2374 1221 -2364
rect 1169 -2544 1221 -2534
rect 1365 -2374 1417 -2364
rect 1365 -2544 1417 -2534
rect 1561 -2374 1613 -2364
rect 1561 -2544 1613 -2534
rect 1757 -2374 1809 -2364
rect 1757 -2544 1809 -2534
rect 1953 -2374 2005 -2364
rect 1953 -2544 2005 -2534
rect 2149 -2374 2201 -2364
rect 2149 -2544 2201 -2534
rect 2345 -2374 2397 -2364
rect 2345 -2544 2397 -2534
rect 2541 -2374 2593 -2364
rect 2541 -2544 2593 -2534
rect 2737 -2374 2789 -2364
rect 2737 -2544 2789 -2534
rect 2933 -2374 2985 -2364
rect 2933 -2544 2985 -2534
rect 679 -2614 731 -2604
rect 679 -2784 731 -2774
rect 875 -2614 927 -2604
rect 875 -2784 927 -2774
rect 1071 -2614 1123 -2604
rect 1071 -2784 1123 -2774
rect 1267 -2614 1319 -2604
rect 1267 -2784 1319 -2774
rect 1463 -2614 1515 -2604
rect 1463 -2784 1515 -2774
rect 1659 -2614 1711 -2604
rect 1659 -2784 1711 -2774
rect 1855 -2614 1907 -2604
rect 1855 -2784 1907 -2774
rect 2051 -2614 2103 -2604
rect 2051 -2784 2103 -2774
rect 2247 -2614 2299 -2604
rect 2247 -2784 2299 -2774
rect 2443 -2614 2495 -2604
rect 2443 -2784 2495 -2774
rect 2639 -2614 2691 -2604
rect 2639 -2784 2691 -2774
rect 2835 -2614 2887 -2604
rect 2835 -2784 2887 -2774
rect 3031 -2614 3083 -2604
rect 3031 -2784 3083 -2774
use sky130_fd_pr__nfet_01v8_lvt_ZRA4RB  sky130_fd_pr__nfet_01v8_lvt_ZRA4RB_0
timestamp 1646921651
transform 1 0 1832 0 1 -2265
box -1392 -719 1392 719
use sky130_fd_pr__nfet_01v8_lvt_ZRA4RB  sky130_fd_pr__nfet_01v8_lvt_ZRA4RB_1
timestamp 1646921651
transform 1 0 1832 0 1 -821
box -1392 -719 1392 719
use sky130_fd_pr__pfet_01v8_NZHYX4  sky130_fd_pr__pfet_01v8_NZHYX4_1
timestamp 1646921651
transform 1 0 1342 0 1 637
box -902 -737 902 737
use sky130_fd_pr__pfet_01v8_NZHYX4  sky130_fd_pr__pfet_01v8_NZHYX4_2
timestamp 1646921651
transform 1 0 3140 0 1 637
box -902 -737 902 737
<< end >>
