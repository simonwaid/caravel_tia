magic
tech sky130A
magscale 1 2
timestamp 1646921651
<< error_p >>
rect -461 981 -403 987
rect -269 981 -211 987
rect -77 981 -19 987
rect 115 981 173 987
rect 307 981 365 987
rect -461 947 -449 981
rect -269 947 -257 981
rect -77 947 -65 981
rect 115 947 127 981
rect 307 947 319 981
rect -461 941 -403 947
rect -269 941 -211 947
rect -77 941 -19 947
rect 115 941 173 947
rect 307 941 365 947
rect -365 71 -307 77
rect -173 71 -115 77
rect 19 71 77 77
rect 211 71 269 77
rect 403 71 461 77
rect -365 37 -353 71
rect -173 37 -161 71
rect 19 37 31 71
rect 211 37 223 71
rect 403 37 415 71
rect -365 31 -307 37
rect -173 31 -115 37
rect 19 31 77 37
rect 211 31 269 37
rect 403 31 461 37
rect -365 -37 -307 -31
rect -173 -37 -115 -31
rect 19 -37 77 -31
rect 211 -37 269 -31
rect 403 -37 461 -31
rect -365 -71 -353 -37
rect -173 -71 -161 -37
rect 19 -71 31 -37
rect 211 -71 223 -37
rect 403 -71 415 -37
rect -365 -77 -307 -71
rect -173 -77 -115 -71
rect 19 -77 77 -71
rect 211 -77 269 -71
rect 403 -77 461 -71
rect -461 -947 -403 -941
rect -269 -947 -211 -941
rect -77 -947 -19 -941
rect 115 -947 173 -941
rect 307 -947 365 -941
rect -461 -981 -449 -947
rect -269 -981 -257 -947
rect -77 -981 -65 -947
rect 115 -981 127 -947
rect 307 -981 319 -947
rect -461 -987 -403 -981
rect -269 -987 -211 -981
rect -77 -987 -19 -981
rect 115 -987 173 -981
rect 307 -987 365 -981
<< pwell >>
rect -647 -1119 647 1119
<< nmoslvt >>
rect -447 109 -417 909
rect -351 109 -321 909
rect -255 109 -225 909
rect -159 109 -129 909
rect -63 109 -33 909
rect 33 109 63 909
rect 129 109 159 909
rect 225 109 255 909
rect 321 109 351 909
rect 417 109 447 909
rect -447 -909 -417 -109
rect -351 -909 -321 -109
rect -255 -909 -225 -109
rect -159 -909 -129 -109
rect -63 -909 -33 -109
rect 33 -909 63 -109
rect 129 -909 159 -109
rect 225 -909 255 -109
rect 321 -909 351 -109
rect 417 -909 447 -109
<< ndiff >>
rect -509 897 -447 909
rect -509 121 -497 897
rect -463 121 -447 897
rect -509 109 -447 121
rect -417 897 -351 909
rect -417 121 -401 897
rect -367 121 -351 897
rect -417 109 -351 121
rect -321 897 -255 909
rect -321 121 -305 897
rect -271 121 -255 897
rect -321 109 -255 121
rect -225 897 -159 909
rect -225 121 -209 897
rect -175 121 -159 897
rect -225 109 -159 121
rect -129 897 -63 909
rect -129 121 -113 897
rect -79 121 -63 897
rect -129 109 -63 121
rect -33 897 33 909
rect -33 121 -17 897
rect 17 121 33 897
rect -33 109 33 121
rect 63 897 129 909
rect 63 121 79 897
rect 113 121 129 897
rect 63 109 129 121
rect 159 897 225 909
rect 159 121 175 897
rect 209 121 225 897
rect 159 109 225 121
rect 255 897 321 909
rect 255 121 271 897
rect 305 121 321 897
rect 255 109 321 121
rect 351 897 417 909
rect 351 121 367 897
rect 401 121 417 897
rect 351 109 417 121
rect 447 897 509 909
rect 447 121 463 897
rect 497 121 509 897
rect 447 109 509 121
rect -509 -121 -447 -109
rect -509 -897 -497 -121
rect -463 -897 -447 -121
rect -509 -909 -447 -897
rect -417 -121 -351 -109
rect -417 -897 -401 -121
rect -367 -897 -351 -121
rect -417 -909 -351 -897
rect -321 -121 -255 -109
rect -321 -897 -305 -121
rect -271 -897 -255 -121
rect -321 -909 -255 -897
rect -225 -121 -159 -109
rect -225 -897 -209 -121
rect -175 -897 -159 -121
rect -225 -909 -159 -897
rect -129 -121 -63 -109
rect -129 -897 -113 -121
rect -79 -897 -63 -121
rect -129 -909 -63 -897
rect -33 -121 33 -109
rect -33 -897 -17 -121
rect 17 -897 33 -121
rect -33 -909 33 -897
rect 63 -121 129 -109
rect 63 -897 79 -121
rect 113 -897 129 -121
rect 63 -909 129 -897
rect 159 -121 225 -109
rect 159 -897 175 -121
rect 209 -897 225 -121
rect 159 -909 225 -897
rect 255 -121 321 -109
rect 255 -897 271 -121
rect 305 -897 321 -121
rect 255 -909 321 -897
rect 351 -121 417 -109
rect 351 -897 367 -121
rect 401 -897 417 -121
rect 351 -909 417 -897
rect 447 -121 509 -109
rect 447 -897 463 -121
rect 497 -897 509 -121
rect 447 -909 509 -897
<< ndiffc >>
rect -497 121 -463 897
rect -401 121 -367 897
rect -305 121 -271 897
rect -209 121 -175 897
rect -113 121 -79 897
rect -17 121 17 897
rect 79 121 113 897
rect 175 121 209 897
rect 271 121 305 897
rect 367 121 401 897
rect 463 121 497 897
rect -497 -897 -463 -121
rect -401 -897 -367 -121
rect -305 -897 -271 -121
rect -209 -897 -175 -121
rect -113 -897 -79 -121
rect -17 -897 17 -121
rect 79 -897 113 -121
rect 175 -897 209 -121
rect 271 -897 305 -121
rect 367 -897 401 -121
rect 463 -897 497 -121
<< psubdiff >>
rect -611 1049 -515 1083
rect 515 1049 611 1083
rect -611 987 -577 1049
rect 577 987 611 1049
rect -611 -1049 -577 -987
rect 577 -1049 611 -987
rect -611 -1083 -515 -1049
rect 515 -1083 611 -1049
<< psubdiffcont >>
rect -515 1049 515 1083
rect -611 -987 -577 987
rect 577 -987 611 987
rect -515 -1083 515 -1049
<< poly >>
rect -465 981 -399 997
rect -465 947 -449 981
rect -415 947 -399 981
rect -465 931 -399 947
rect -273 981 -207 997
rect -273 947 -257 981
rect -223 947 -207 981
rect -447 909 -417 931
rect -351 909 -321 935
rect -273 931 -207 947
rect -81 981 -15 997
rect -81 947 -65 981
rect -31 947 -15 981
rect -255 909 -225 931
rect -159 909 -129 935
rect -81 931 -15 947
rect 111 981 177 997
rect 111 947 127 981
rect 161 947 177 981
rect -63 909 -33 931
rect 33 909 63 935
rect 111 931 177 947
rect 303 981 369 997
rect 303 947 319 981
rect 353 947 369 981
rect 129 909 159 931
rect 225 909 255 935
rect 303 931 369 947
rect 321 909 351 931
rect 417 909 447 935
rect -447 83 -417 109
rect -351 87 -321 109
rect -369 71 -303 87
rect -255 83 -225 109
rect -159 87 -129 109
rect -369 37 -353 71
rect -319 37 -303 71
rect -369 21 -303 37
rect -177 71 -111 87
rect -63 83 -33 109
rect 33 87 63 109
rect -177 37 -161 71
rect -127 37 -111 71
rect -177 21 -111 37
rect 15 71 81 87
rect 129 83 159 109
rect 225 87 255 109
rect 15 37 31 71
rect 65 37 81 71
rect 15 21 81 37
rect 207 71 273 87
rect 321 83 351 109
rect 417 87 447 109
rect 207 37 223 71
rect 257 37 273 71
rect 207 21 273 37
rect 399 71 465 87
rect 399 37 415 71
rect 449 37 465 71
rect 399 21 465 37
rect -369 -37 -303 -21
rect -369 -71 -353 -37
rect -319 -71 -303 -37
rect -447 -109 -417 -83
rect -369 -87 -303 -71
rect -177 -37 -111 -21
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect -351 -109 -321 -87
rect -255 -109 -225 -83
rect -177 -87 -111 -71
rect 15 -37 81 -21
rect 15 -71 31 -37
rect 65 -71 81 -37
rect -159 -109 -129 -87
rect -63 -109 -33 -83
rect 15 -87 81 -71
rect 207 -37 273 -21
rect 207 -71 223 -37
rect 257 -71 273 -37
rect 33 -109 63 -87
rect 129 -109 159 -83
rect 207 -87 273 -71
rect 399 -37 465 -21
rect 399 -71 415 -37
rect 449 -71 465 -37
rect 225 -109 255 -87
rect 321 -109 351 -83
rect 399 -87 465 -71
rect 417 -109 447 -87
rect -447 -931 -417 -909
rect -465 -947 -399 -931
rect -351 -935 -321 -909
rect -255 -931 -225 -909
rect -465 -981 -449 -947
rect -415 -981 -399 -947
rect -465 -997 -399 -981
rect -273 -947 -207 -931
rect -159 -935 -129 -909
rect -63 -931 -33 -909
rect -273 -981 -257 -947
rect -223 -981 -207 -947
rect -273 -997 -207 -981
rect -81 -947 -15 -931
rect 33 -935 63 -909
rect 129 -931 159 -909
rect -81 -981 -65 -947
rect -31 -981 -15 -947
rect -81 -997 -15 -981
rect 111 -947 177 -931
rect 225 -935 255 -909
rect 321 -931 351 -909
rect 111 -981 127 -947
rect 161 -981 177 -947
rect 111 -997 177 -981
rect 303 -947 369 -931
rect 417 -935 447 -909
rect 303 -981 319 -947
rect 353 -981 369 -947
rect 303 -997 369 -981
<< polycont >>
rect -449 947 -415 981
rect -257 947 -223 981
rect -65 947 -31 981
rect 127 947 161 981
rect 319 947 353 981
rect -353 37 -319 71
rect -161 37 -127 71
rect 31 37 65 71
rect 223 37 257 71
rect 415 37 449 71
rect -353 -71 -319 -37
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect 223 -71 257 -37
rect 415 -71 449 -37
rect -449 -981 -415 -947
rect -257 -981 -223 -947
rect -65 -981 -31 -947
rect 127 -981 161 -947
rect 319 -981 353 -947
<< locali >>
rect -611 1049 -515 1083
rect 515 1049 611 1083
rect -611 987 -577 1049
rect 577 987 611 1049
rect -465 947 -449 981
rect -415 947 -399 981
rect -273 947 -257 981
rect -223 947 -207 981
rect -81 947 -65 981
rect -31 947 -15 981
rect 111 947 127 981
rect 161 947 177 981
rect 303 947 319 981
rect 353 947 369 981
rect -497 897 -463 913
rect -497 105 -463 121
rect -401 897 -367 913
rect -401 105 -367 121
rect -305 897 -271 913
rect -305 105 -271 121
rect -209 897 -175 913
rect -209 105 -175 121
rect -113 897 -79 913
rect -113 105 -79 121
rect -17 897 17 913
rect -17 105 17 121
rect 79 897 113 913
rect 79 105 113 121
rect 175 897 209 913
rect 175 105 209 121
rect 271 897 305 913
rect 271 105 305 121
rect 367 897 401 913
rect 367 105 401 121
rect 463 897 497 913
rect 463 105 497 121
rect -369 37 -353 71
rect -319 37 -303 71
rect -177 37 -161 71
rect -127 37 -111 71
rect 15 37 31 71
rect 65 37 81 71
rect 207 37 223 71
rect 257 37 273 71
rect 399 37 415 71
rect 449 37 465 71
rect -369 -71 -353 -37
rect -319 -71 -303 -37
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect 15 -71 31 -37
rect 65 -71 81 -37
rect 207 -71 223 -37
rect 257 -71 273 -37
rect 399 -71 415 -37
rect 449 -71 465 -37
rect -497 -121 -463 -105
rect -497 -913 -463 -897
rect -401 -121 -367 -105
rect -401 -913 -367 -897
rect -305 -121 -271 -105
rect -305 -913 -271 -897
rect -209 -121 -175 -105
rect -209 -913 -175 -897
rect -113 -121 -79 -105
rect -113 -913 -79 -897
rect -17 -121 17 -105
rect -17 -913 17 -897
rect 79 -121 113 -105
rect 79 -913 113 -897
rect 175 -121 209 -105
rect 175 -913 209 -897
rect 271 -121 305 -105
rect 271 -913 305 -897
rect 367 -121 401 -105
rect 367 -913 401 -897
rect 463 -121 497 -105
rect 463 -913 497 -897
rect -465 -981 -449 -947
rect -415 -981 -399 -947
rect -273 -981 -257 -947
rect -223 -981 -207 -947
rect -81 -981 -65 -947
rect -31 -981 -15 -947
rect 111 -981 127 -947
rect 161 -981 177 -947
rect 303 -981 319 -947
rect 353 -981 369 -947
rect -611 -1049 -577 -987
rect 577 -1049 611 -987
rect -611 -1083 -515 -1049
rect 515 -1083 611 -1049
<< viali >>
rect -449 947 -415 981
rect -257 947 -223 981
rect -65 947 -31 981
rect 127 947 161 981
rect 319 947 353 981
rect -497 121 -463 897
rect -401 121 -367 897
rect -305 121 -271 897
rect -209 121 -175 897
rect -113 121 -79 897
rect -17 121 17 897
rect 79 121 113 897
rect 175 121 209 897
rect 271 121 305 897
rect 367 121 401 897
rect 463 121 497 897
rect -353 37 -319 71
rect -161 37 -127 71
rect 31 37 65 71
rect 223 37 257 71
rect 415 37 449 71
rect -353 -71 -319 -37
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect 223 -71 257 -37
rect 415 -71 449 -37
rect -497 -897 -463 -121
rect -401 -897 -367 -121
rect -305 -897 -271 -121
rect -209 -897 -175 -121
rect -113 -897 -79 -121
rect -17 -897 17 -121
rect 79 -897 113 -121
rect 175 -897 209 -121
rect 271 -897 305 -121
rect 367 -897 401 -121
rect 463 -897 497 -121
rect -449 -981 -415 -947
rect -257 -981 -223 -947
rect -65 -981 -31 -947
rect 127 -981 161 -947
rect 319 -981 353 -947
<< metal1 >>
rect -461 981 -403 987
rect -461 947 -449 981
rect -415 947 -403 981
rect -461 941 -403 947
rect -269 981 -211 987
rect -269 947 -257 981
rect -223 947 -211 981
rect -269 941 -211 947
rect -77 981 -19 987
rect -77 947 -65 981
rect -31 947 -19 981
rect -77 941 -19 947
rect 115 981 173 987
rect 115 947 127 981
rect 161 947 173 981
rect 115 941 173 947
rect 307 981 365 987
rect 307 947 319 981
rect 353 947 365 981
rect 307 941 365 947
rect -503 897 -457 909
rect -503 121 -497 897
rect -463 121 -457 897
rect -503 109 -457 121
rect -407 897 -361 909
rect -407 121 -401 897
rect -367 121 -361 897
rect -407 109 -361 121
rect -311 897 -265 909
rect -311 121 -305 897
rect -271 121 -265 897
rect -311 109 -265 121
rect -215 897 -169 909
rect -215 121 -209 897
rect -175 121 -169 897
rect -215 109 -169 121
rect -119 897 -73 909
rect -119 121 -113 897
rect -79 121 -73 897
rect -119 109 -73 121
rect -23 897 23 909
rect -23 121 -17 897
rect 17 121 23 897
rect -23 109 23 121
rect 73 897 119 909
rect 73 121 79 897
rect 113 121 119 897
rect 73 109 119 121
rect 169 897 215 909
rect 169 121 175 897
rect 209 121 215 897
rect 169 109 215 121
rect 265 897 311 909
rect 265 121 271 897
rect 305 121 311 897
rect 265 109 311 121
rect 361 897 407 909
rect 361 121 367 897
rect 401 121 407 897
rect 361 109 407 121
rect 457 897 503 909
rect 457 121 463 897
rect 497 121 503 897
rect 457 109 503 121
rect -365 71 -307 77
rect -365 37 -353 71
rect -319 37 -307 71
rect -365 31 -307 37
rect -173 71 -115 77
rect -173 37 -161 71
rect -127 37 -115 71
rect -173 31 -115 37
rect 19 71 77 77
rect 19 37 31 71
rect 65 37 77 71
rect 19 31 77 37
rect 211 71 269 77
rect 211 37 223 71
rect 257 37 269 71
rect 211 31 269 37
rect 403 71 461 77
rect 403 37 415 71
rect 449 37 461 71
rect 403 31 461 37
rect -365 -37 -307 -31
rect -365 -71 -353 -37
rect -319 -71 -307 -37
rect -365 -77 -307 -71
rect -173 -37 -115 -31
rect -173 -71 -161 -37
rect -127 -71 -115 -37
rect -173 -77 -115 -71
rect 19 -37 77 -31
rect 19 -71 31 -37
rect 65 -71 77 -37
rect 19 -77 77 -71
rect 211 -37 269 -31
rect 211 -71 223 -37
rect 257 -71 269 -37
rect 211 -77 269 -71
rect 403 -37 461 -31
rect 403 -71 415 -37
rect 449 -71 461 -37
rect 403 -77 461 -71
rect -503 -121 -457 -109
rect -503 -897 -497 -121
rect -463 -897 -457 -121
rect -503 -909 -457 -897
rect -407 -121 -361 -109
rect -407 -897 -401 -121
rect -367 -897 -361 -121
rect -407 -909 -361 -897
rect -311 -121 -265 -109
rect -311 -897 -305 -121
rect -271 -897 -265 -121
rect -311 -909 -265 -897
rect -215 -121 -169 -109
rect -215 -897 -209 -121
rect -175 -897 -169 -121
rect -215 -909 -169 -897
rect -119 -121 -73 -109
rect -119 -897 -113 -121
rect -79 -897 -73 -121
rect -119 -909 -73 -897
rect -23 -121 23 -109
rect -23 -897 -17 -121
rect 17 -897 23 -121
rect -23 -909 23 -897
rect 73 -121 119 -109
rect 73 -897 79 -121
rect 113 -897 119 -121
rect 73 -909 119 -897
rect 169 -121 215 -109
rect 169 -897 175 -121
rect 209 -897 215 -121
rect 169 -909 215 -897
rect 265 -121 311 -109
rect 265 -897 271 -121
rect 305 -897 311 -121
rect 265 -909 311 -897
rect 361 -121 407 -109
rect 361 -897 367 -121
rect 401 -897 407 -121
rect 361 -909 407 -897
rect 457 -121 503 -109
rect 457 -897 463 -121
rect 497 -897 503 -121
rect 457 -909 503 -897
rect -461 -947 -403 -941
rect -461 -981 -449 -947
rect -415 -981 -403 -947
rect -461 -987 -403 -981
rect -269 -947 -211 -941
rect -269 -981 -257 -947
rect -223 -981 -211 -947
rect -269 -987 -211 -981
rect -77 -947 -19 -941
rect -77 -981 -65 -947
rect -31 -981 -19 -947
rect -77 -987 -19 -981
rect 115 -947 173 -941
rect 115 -981 127 -947
rect 161 -981 173 -947
rect 115 -987 173 -981
rect 307 -947 365 -941
rect 307 -981 319 -947
rect 353 -981 365 -947
rect 307 -987 365 -981
<< properties >>
string FIXED_BBOX -594 -1066 594 1066
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 4 l 0.150 m 2 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
