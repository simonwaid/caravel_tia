magic
tech sky130A
timestamp 1646682533
<< nwell >>
rect -2351 269 281 507
<< pwell >>
rect -2420 507 350 576
rect -2420 269 -2351 507
rect 281 269 350 507
rect -2420 200 350 269
rect -2350 -40 282 198
<< psubdiff >>
rect -2402 541 -2354 558
rect 284 541 332 558
rect -2402 510 -2385 541
rect 315 510 332 541
rect -2402 235 -2385 266
rect 315 235 332 266
rect -2402 218 -2354 235
rect 284 218 332 235
rect -2332 163 -2284 180
rect -2178 163 -2130 180
rect -2332 132 -2315 163
rect -2147 132 -2130 163
rect -2332 -5 -2315 26
rect -2147 -5 -2130 26
rect -2332 -22 -2284 -5
rect -2178 -22 -2130 -5
rect -2066 163 -2018 180
rect -1912 163 -1864 180
rect -2066 132 -2049 163
rect -1881 132 -1864 163
rect -2066 -5 -2049 26
rect -1881 -5 -1864 26
rect -2066 -22 -2018 -5
rect -1912 -22 -1864 -5
rect -1800 163 -1752 180
rect -1646 163 -1598 180
rect -1800 132 -1783 163
rect -1615 132 -1598 163
rect -1800 -5 -1783 26
rect -1615 -5 -1598 26
rect -1800 -22 -1752 -5
rect -1646 -22 -1598 -5
rect -1534 163 -1486 180
rect -1380 163 -1332 180
rect -1534 132 -1517 163
rect -1349 132 -1332 163
rect -1534 -5 -1517 26
rect -1349 -5 -1332 26
rect -1534 -22 -1486 -5
rect -1380 -22 -1332 -5
rect -1268 163 -1220 180
rect -1114 163 -1066 180
rect -1268 132 -1251 163
rect -1083 132 -1066 163
rect -1268 -5 -1251 26
rect -1083 -5 -1066 26
rect -1268 -22 -1220 -5
rect -1114 -22 -1066 -5
rect -1002 163 -954 180
rect -848 163 -800 180
rect -1002 132 -985 163
rect -817 132 -800 163
rect -1002 -5 -985 26
rect -817 -5 -800 26
rect -1002 -22 -954 -5
rect -848 -22 -800 -5
rect -736 163 -688 180
rect -582 163 -534 180
rect -736 132 -719 163
rect -551 132 -534 163
rect -736 -5 -719 26
rect -551 -5 -534 26
rect -736 -22 -688 -5
rect -582 -22 -534 -5
rect -470 163 -422 180
rect -316 163 -268 180
rect -470 132 -453 163
rect -285 132 -268 163
rect -470 -5 -453 26
rect -285 -5 -268 26
rect -470 -22 -422 -5
rect -316 -22 -268 -5
rect -204 163 -156 180
rect -50 163 -2 180
rect -204 132 -187 163
rect -19 132 -2 163
rect -204 -5 -187 26
rect -19 -5 -2 26
rect -204 -22 -156 -5
rect -50 -22 -2 -5
rect 62 163 110 180
rect 216 163 264 180
rect 62 132 79 163
rect 247 132 264 163
rect 62 -5 79 26
rect 247 -5 264 26
rect 62 -22 110 -5
rect 216 -22 264 -5
<< nsubdiff >>
rect -2333 472 -2285 489
rect -2179 472 -2131 489
rect -2333 441 -2316 472
rect -2148 441 -2131 472
rect -2333 304 -2316 335
rect -2148 304 -2131 335
rect -2333 287 -2285 304
rect -2179 287 -2131 304
rect -2067 472 -2019 489
rect -1913 472 -1865 489
rect -2067 441 -2050 472
rect -1882 441 -1865 472
rect -2067 304 -2050 335
rect -1882 304 -1865 335
rect -2067 287 -2019 304
rect -1913 287 -1865 304
rect -1801 472 -1753 489
rect -1647 472 -1599 489
rect -1801 441 -1784 472
rect -1616 441 -1599 472
rect -1801 304 -1784 335
rect -1616 304 -1599 335
rect -1801 287 -1753 304
rect -1647 287 -1599 304
rect -1535 472 -1487 489
rect -1381 472 -1333 489
rect -1535 441 -1518 472
rect -1350 441 -1333 472
rect -1535 304 -1518 335
rect -1350 304 -1333 335
rect -1535 287 -1487 304
rect -1381 287 -1333 304
rect -1269 472 -1221 489
rect -1115 472 -1067 489
rect -1269 441 -1252 472
rect -1084 441 -1067 472
rect -1269 304 -1252 335
rect -1084 304 -1067 335
rect -1269 287 -1221 304
rect -1115 287 -1067 304
rect -1003 472 -955 489
rect -849 472 -801 489
rect -1003 441 -986 472
rect -818 441 -801 472
rect -1003 304 -986 335
rect -818 304 -801 335
rect -1003 287 -955 304
rect -849 287 -801 304
rect -737 472 -689 489
rect -583 472 -535 489
rect -737 441 -720 472
rect -552 441 -535 472
rect -737 304 -720 335
rect -552 304 -535 335
rect -737 287 -689 304
rect -583 287 -535 304
rect -471 472 -423 489
rect -317 472 -269 489
rect -471 441 -454 472
rect -286 441 -269 472
rect -471 304 -454 335
rect -286 304 -269 335
rect -471 287 -423 304
rect -317 287 -269 304
rect -205 472 -157 489
rect -51 472 -3 489
rect -205 441 -188 472
rect -20 441 -3 472
rect -205 304 -188 335
rect -20 304 -3 335
rect -205 287 -157 304
rect -51 287 -3 304
rect 61 472 109 489
rect 215 472 263 489
rect 61 441 78 472
rect 246 441 263 472
rect 61 304 78 335
rect 246 304 263 335
rect 61 287 109 304
rect 215 287 263 304
<< psubdiffcont >>
rect -2354 541 284 558
rect -2402 266 -2385 510
rect 315 266 332 510
rect -2354 218 284 235
rect -2284 163 -2178 180
rect -2332 26 -2315 132
rect -2147 26 -2130 132
rect -2284 -22 -2178 -5
rect -2018 163 -1912 180
rect -2066 26 -2049 132
rect -1881 26 -1864 132
rect -2018 -22 -1912 -5
rect -1752 163 -1646 180
rect -1800 26 -1783 132
rect -1615 26 -1598 132
rect -1752 -22 -1646 -5
rect -1486 163 -1380 180
rect -1534 26 -1517 132
rect -1349 26 -1332 132
rect -1486 -22 -1380 -5
rect -1220 163 -1114 180
rect -1268 26 -1251 132
rect -1083 26 -1066 132
rect -1220 -22 -1114 -5
rect -954 163 -848 180
rect -1002 26 -985 132
rect -817 26 -800 132
rect -954 -22 -848 -5
rect -688 163 -582 180
rect -736 26 -719 132
rect -551 26 -534 132
rect -688 -22 -582 -5
rect -422 163 -316 180
rect -470 26 -453 132
rect -285 26 -268 132
rect -422 -22 -316 -5
rect -156 163 -50 180
rect -204 26 -187 132
rect -19 26 -2 132
rect -156 -22 -50 -5
rect 110 163 216 180
rect 62 26 79 132
rect 247 26 264 132
rect 110 -22 216 -5
<< nsubdiffcont >>
rect -2285 472 -2179 489
rect -2333 335 -2316 441
rect -2148 335 -2131 441
rect -2285 287 -2179 304
rect -2019 472 -1913 489
rect -2067 335 -2050 441
rect -1882 335 -1865 441
rect -2019 287 -1913 304
rect -1753 472 -1647 489
rect -1801 335 -1784 441
rect -1616 335 -1599 441
rect -1753 287 -1647 304
rect -1487 472 -1381 489
rect -1535 335 -1518 441
rect -1350 335 -1333 441
rect -1487 287 -1381 304
rect -1221 472 -1115 489
rect -1269 335 -1252 441
rect -1084 335 -1067 441
rect -1221 287 -1115 304
rect -955 472 -849 489
rect -1003 335 -986 441
rect -818 335 -801 441
rect -955 287 -849 304
rect -689 472 -583 489
rect -737 335 -720 441
rect -552 335 -535 441
rect -689 287 -583 304
rect -423 472 -317 489
rect -471 335 -454 441
rect -286 335 -269 441
rect -423 287 -317 304
rect -157 472 -51 489
rect -205 335 -188 441
rect -20 335 -3 441
rect -157 287 -51 304
rect 109 472 215 489
rect 61 335 78 441
rect 246 335 263 441
rect 109 287 215 304
<< pdiode >>
rect -2282 432 -2182 438
rect -2282 344 -2276 432
rect -2188 344 -2182 432
rect -2282 338 -2182 344
rect -2016 432 -1916 438
rect -2016 344 -2010 432
rect -1922 344 -1916 432
rect -2016 338 -1916 344
rect -1750 432 -1650 438
rect -1750 344 -1744 432
rect -1656 344 -1650 432
rect -1750 338 -1650 344
rect -1484 432 -1384 438
rect -1484 344 -1478 432
rect -1390 344 -1384 432
rect -1484 338 -1384 344
rect -1218 432 -1118 438
rect -1218 344 -1212 432
rect -1124 344 -1118 432
rect -1218 338 -1118 344
rect -952 432 -852 438
rect -952 344 -946 432
rect -858 344 -852 432
rect -952 338 -852 344
rect -686 432 -586 438
rect -686 344 -680 432
rect -592 344 -586 432
rect -686 338 -586 344
rect -420 432 -320 438
rect -420 344 -414 432
rect -326 344 -320 432
rect -420 338 -320 344
rect -154 432 -54 438
rect -154 344 -148 432
rect -60 344 -54 432
rect -154 338 -54 344
rect 112 432 212 438
rect 112 344 118 432
rect 206 344 212 432
rect 112 338 212 344
<< ndiode >>
rect -2281 123 -2181 129
rect -2281 35 -2275 123
rect -2187 35 -2181 123
rect -2281 29 -2181 35
rect -2015 123 -1915 129
rect -2015 35 -2009 123
rect -1921 35 -1915 123
rect -2015 29 -1915 35
rect -1749 123 -1649 129
rect -1749 35 -1743 123
rect -1655 35 -1649 123
rect -1749 29 -1649 35
rect -1483 123 -1383 129
rect -1483 35 -1477 123
rect -1389 35 -1383 123
rect -1483 29 -1383 35
rect -1217 123 -1117 129
rect -1217 35 -1211 123
rect -1123 35 -1117 123
rect -1217 29 -1117 35
rect -951 123 -851 129
rect -951 35 -945 123
rect -857 35 -851 123
rect -951 29 -851 35
rect -685 123 -585 129
rect -685 35 -679 123
rect -591 35 -585 123
rect -685 29 -585 35
rect -419 123 -319 129
rect -419 35 -413 123
rect -325 35 -319 123
rect -419 29 -319 35
rect -153 123 -53 129
rect -153 35 -147 123
rect -59 35 -53 123
rect -153 29 -53 35
rect 113 123 213 129
rect 113 35 119 123
rect 207 35 213 123
rect 113 29 213 35
<< pdiodec >>
rect -2276 344 -2188 432
rect -2010 344 -1922 432
rect -1744 344 -1656 432
rect -1478 344 -1390 432
rect -1212 344 -1124 432
rect -946 344 -858 432
rect -680 344 -592 432
rect -414 344 -326 432
rect -148 344 -60 432
rect 118 344 206 432
<< ndiodec >>
rect -2275 35 -2187 123
rect -2009 35 -1921 123
rect -1743 35 -1655 123
rect -1477 35 -1389 123
rect -1211 35 -1123 123
rect -945 35 -857 123
rect -679 35 -591 123
rect -413 35 -325 123
rect -147 35 -59 123
rect 119 35 207 123
<< locali >>
rect -2420 558 350 575
rect -2420 541 -2354 558
rect 284 541 350 558
rect -2420 510 -2385 541
rect -2420 266 -2402 510
rect 315 510 350 541
rect -2350 489 280 505
rect -2350 472 -2285 489
rect -2179 472 -2019 489
rect -1913 472 -1753 489
rect -1647 472 -1487 489
rect -1381 472 -1221 489
rect -1115 472 -955 489
rect -849 472 -689 489
rect -583 472 -423 489
rect -317 472 -157 489
rect -51 472 109 489
rect 215 472 280 489
rect -2350 441 -2316 472
rect -2350 335 -2333 441
rect -2148 441 -2050 472
rect -2284 344 -2276 432
rect -2188 344 -2180 432
rect -2350 304 -2316 335
rect -2131 335 -2067 441
rect -1882 441 -1784 472
rect -2018 344 -2010 432
rect -1922 344 -1914 432
rect -2148 304 -2050 335
rect -1865 335 -1801 441
rect -1616 441 -1518 472
rect -1752 344 -1744 432
rect -1656 344 -1648 432
rect -1882 304 -1784 335
rect -1599 335 -1535 441
rect -1350 441 -1252 472
rect -1486 344 -1478 432
rect -1390 344 -1382 432
rect -1616 304 -1518 335
rect -1333 335 -1269 441
rect -1084 441 -986 472
rect -1220 344 -1212 432
rect -1124 344 -1116 432
rect -1350 304 -1252 335
rect -1067 335 -1003 441
rect -818 441 -720 472
rect -954 344 -946 432
rect -858 344 -850 432
rect -1084 304 -986 335
rect -801 335 -737 441
rect -552 441 -454 472
rect -688 344 -680 432
rect -592 344 -584 432
rect -818 304 -720 335
rect -535 335 -471 441
rect -286 441 -188 472
rect -422 344 -414 432
rect -326 344 -318 432
rect -552 304 -454 335
rect -269 335 -205 441
rect -20 441 78 472
rect -156 344 -148 432
rect -60 344 -52 432
rect -286 304 -188 335
rect -3 335 61 441
rect 246 441 280 472
rect 110 344 118 432
rect 206 344 214 432
rect -20 304 78 335
rect 263 335 280 441
rect 246 304 280 335
rect -2350 287 -2285 304
rect -2179 287 -2019 304
rect -1913 287 -1753 304
rect -1647 287 -1487 304
rect -1381 287 -1221 304
rect -1115 287 -955 304
rect -849 287 -689 304
rect -583 287 -423 304
rect -317 287 -157 304
rect -51 287 109 304
rect 215 287 280 304
rect -2350 270 280 287
rect -2420 235 -2385 266
rect 332 266 350 510
rect 315 235 350 266
rect -2420 218 -2354 235
rect 284 218 350 235
rect -2420 180 350 218
rect -2420 163 -2284 180
rect -2178 163 -2018 180
rect -1912 163 -1752 180
rect -1646 163 -1486 180
rect -1380 163 -1220 180
rect -1114 163 -954 180
rect -848 163 -688 180
rect -582 163 -422 180
rect -316 163 -156 180
rect -50 163 110 180
rect 216 163 350 180
rect -2420 132 -2315 163
rect -2420 26 -2332 132
rect -2147 132 -2049 163
rect -2283 35 -2275 123
rect -2187 35 -2179 123
rect -2420 -5 -2315 26
rect -2130 26 -2066 132
rect -1881 132 -1783 163
rect -2017 35 -2009 123
rect -1921 35 -1913 123
rect -2147 -5 -2049 26
rect -1864 26 -1800 132
rect -1615 132 -1517 163
rect -1751 35 -1743 123
rect -1655 35 -1647 123
rect -1881 -5 -1783 26
rect -1598 26 -1534 132
rect -1349 132 -1251 163
rect -1485 35 -1477 123
rect -1389 35 -1381 123
rect -1615 -5 -1517 26
rect -1332 26 -1268 132
rect -1083 132 -985 163
rect -1219 35 -1211 123
rect -1123 35 -1115 123
rect -1349 -5 -1251 26
rect -1066 26 -1002 132
rect -817 132 -719 163
rect -953 35 -945 123
rect -857 35 -849 123
rect -1083 -5 -985 26
rect -800 26 -736 132
rect -551 132 -453 163
rect -687 35 -679 123
rect -591 35 -583 123
rect -817 -5 -719 26
rect -534 26 -470 132
rect -285 132 -187 163
rect -421 35 -413 123
rect -325 35 -317 123
rect -551 -5 -453 26
rect -268 26 -204 132
rect -19 132 79 163
rect -155 35 -147 123
rect -59 35 -51 123
rect -285 -5 -187 26
rect -2 26 62 132
rect 247 132 350 163
rect 111 35 119 123
rect 207 35 215 123
rect -19 -5 79 26
rect 264 26 350 132
rect 247 -5 350 26
rect -2420 -22 -2284 -5
rect -2178 -22 -2018 -5
rect -1912 -22 -1752 -5
rect -1646 -22 -1486 -5
rect -1380 -22 -1220 -5
rect -1114 -22 -954 -5
rect -848 -22 -688 -5
rect -582 -22 -422 -5
rect -316 -22 -156 -5
rect -50 -22 110 -5
rect 216 -22 350 -5
rect -2420 -45 350 -22
<< viali >>
rect -2276 344 -2188 432
rect -2010 344 -1922 432
rect -1744 344 -1656 432
rect -1478 344 -1390 432
rect -1212 344 -1124 432
rect -946 344 -858 432
rect -680 344 -592 432
rect -414 344 -326 432
rect -148 344 -60 432
rect 118 344 206 432
rect -2275 35 -2187 123
rect -2009 35 -1921 123
rect -1743 35 -1655 123
rect -1477 35 -1389 123
rect -1211 35 -1123 123
rect -945 35 -857 123
rect -679 35 -591 123
rect -413 35 -325 123
rect -147 35 -59 123
rect 119 35 207 123
<< metal1 >>
rect -2282 432 -2182 435
rect -2282 344 -2276 432
rect -2188 344 -2182 432
rect -2282 341 -2182 344
rect -2016 432 -1916 435
rect -2016 344 -2010 432
rect -1922 344 -1916 432
rect -2016 341 -1916 344
rect -1750 432 -1650 435
rect -1750 344 -1744 432
rect -1656 344 -1650 432
rect -1750 341 -1650 344
rect -1484 432 -1384 435
rect -1484 344 -1478 432
rect -1390 344 -1384 432
rect -1484 341 -1384 344
rect -1218 432 -1118 435
rect -1218 344 -1212 432
rect -1124 344 -1118 432
rect -1218 341 -1118 344
rect -952 432 -852 435
rect -952 344 -946 432
rect -858 344 -852 432
rect -952 341 -852 344
rect -686 432 -586 435
rect -686 344 -680 432
rect -592 344 -586 432
rect -686 341 -586 344
rect -420 432 -320 435
rect -420 344 -414 432
rect -326 344 -320 432
rect -420 341 -320 344
rect -154 432 -54 435
rect -154 344 -148 432
rect -60 344 -54 432
rect -154 341 -54 344
rect 112 432 212 435
rect 112 344 118 432
rect 206 344 212 432
rect 112 341 212 344
rect -2281 123 -2181 126
rect -2281 35 -2275 123
rect -2187 35 -2181 123
rect -2281 32 -2181 35
rect -2015 123 -1915 126
rect -2015 35 -2009 123
rect -1921 35 -1915 123
rect -2015 32 -1915 35
rect -1749 123 -1649 126
rect -1749 35 -1743 123
rect -1655 35 -1649 123
rect -1749 32 -1649 35
rect -1483 123 -1383 126
rect -1483 35 -1477 123
rect -1389 35 -1383 123
rect -1483 32 -1383 35
rect -1217 123 -1117 126
rect -1217 35 -1211 123
rect -1123 35 -1117 123
rect -1217 32 -1117 35
rect -951 123 -851 126
rect -951 35 -945 123
rect -857 35 -851 123
rect -951 32 -851 35
rect -685 123 -585 126
rect -685 35 -679 123
rect -591 35 -585 123
rect -685 32 -585 35
rect -419 123 -319 126
rect -419 35 -413 123
rect -325 35 -319 123
rect -419 32 -319 35
rect -153 123 -53 126
rect -153 35 -147 123
rect -59 35 -53 123
rect -153 32 -53 35
rect 113 123 213 126
rect 113 35 119 123
rect 207 35 213 123
rect 113 32 213 35
use sky130_fd_pr__diode_pd2nw_05v5_AEDW7W  sky130_fd_pr__diode_pd2nw_05v5_AEDW7W_0
timestamp 1646653136
transform 1 0 -1035 0 1 388
box -1385 -188 1385 188
use sky130_fd_pr__diode_pw2nd_05v5_Z3EYSA  sky130_fd_pr__diode_pw2nd_05v5_Z3EYSA_0
timestamp 1646653136
transform 1 0 -1034 0 1 79
box -1316 -119 1316 119
<< end >>
