magic
tech sky130A
timestamp 1646921651
<< pwell >>
rect -1656 -305 1656 305
<< nmos >>
rect -1558 -200 -958 200
rect -929 -200 -329 200
rect -300 -200 300 200
rect 329 -200 929 200
rect 958 -200 1558 200
<< ndiff >>
rect -1587 194 -1558 200
rect -1587 -194 -1581 194
rect -1564 -194 -1558 194
rect -1587 -200 -1558 -194
rect -958 194 -929 200
rect -958 -194 -952 194
rect -935 -194 -929 194
rect -958 -200 -929 -194
rect -329 194 -300 200
rect -329 -194 -323 194
rect -306 -194 -300 194
rect -329 -200 -300 -194
rect 300 194 329 200
rect 300 -194 306 194
rect 323 -194 329 194
rect 300 -200 329 -194
rect 929 194 958 200
rect 929 -194 935 194
rect 952 -194 958 194
rect 929 -200 958 -194
rect 1558 194 1587 200
rect 1558 -194 1564 194
rect 1581 -194 1587 194
rect 1558 -200 1587 -194
<< ndiffc >>
rect -1581 -194 -1564 194
rect -952 -194 -935 194
rect -323 -194 -306 194
rect 306 -194 323 194
rect 935 -194 952 194
rect 1564 -194 1581 194
<< psubdiff >>
rect -1638 270 -1590 287
rect 1590 270 1638 287
rect -1638 239 -1621 270
rect 1621 239 1638 270
rect -1638 -270 -1621 -239
rect 1621 -270 1638 -239
rect -1638 -287 -1590 -270
rect 1590 -287 1638 -270
<< psubdiffcont >>
rect -1590 270 1590 287
rect -1638 -239 -1621 239
rect 1621 -239 1638 239
rect -1590 -287 1590 -270
<< poly >>
rect -1558 236 -958 244
rect -1558 219 -1550 236
rect -966 219 -958 236
rect -1558 200 -958 219
rect -929 236 -329 244
rect -929 219 -921 236
rect -337 219 -329 236
rect -929 200 -329 219
rect -300 236 300 244
rect -300 219 -292 236
rect 292 219 300 236
rect -300 200 300 219
rect 329 236 929 244
rect 329 219 337 236
rect 921 219 929 236
rect 329 200 929 219
rect 958 236 1558 244
rect 958 219 966 236
rect 1550 219 1558 236
rect 958 200 1558 219
rect -1558 -219 -958 -200
rect -1558 -236 -1550 -219
rect -966 -236 -958 -219
rect -1558 -244 -958 -236
rect -929 -219 -329 -200
rect -929 -236 -921 -219
rect -337 -236 -329 -219
rect -929 -244 -329 -236
rect -300 -219 300 -200
rect -300 -236 -292 -219
rect 292 -236 300 -219
rect -300 -244 300 -236
rect 329 -219 929 -200
rect 329 -236 337 -219
rect 921 -236 929 -219
rect 329 -244 929 -236
rect 958 -219 1558 -200
rect 958 -236 966 -219
rect 1550 -236 1558 -219
rect 958 -244 1558 -236
<< polycont >>
rect -1550 219 -966 236
rect -921 219 -337 236
rect -292 219 292 236
rect 337 219 921 236
rect 966 219 1550 236
rect -1550 -236 -966 -219
rect -921 -236 -337 -219
rect -292 -236 292 -219
rect 337 -236 921 -219
rect 966 -236 1550 -219
<< locali >>
rect -1638 270 -1590 287
rect 1590 270 1638 287
rect -1638 239 -1621 270
rect 1621 239 1638 270
rect -1558 219 -1550 236
rect -966 219 -958 236
rect -929 219 -921 236
rect -337 219 -329 236
rect -300 219 -292 236
rect 292 219 300 236
rect 329 219 337 236
rect 921 219 929 236
rect 958 219 966 236
rect 1550 219 1558 236
rect -1581 194 -1564 202
rect -1581 -202 -1564 -194
rect -952 194 -935 202
rect -952 -202 -935 -194
rect -323 194 -306 202
rect -323 -202 -306 -194
rect 306 194 323 202
rect 306 -202 323 -194
rect 935 194 952 202
rect 935 -202 952 -194
rect 1564 194 1581 202
rect 1564 -202 1581 -194
rect -1558 -236 -1550 -219
rect -966 -236 -958 -219
rect -929 -236 -921 -219
rect -337 -236 -329 -219
rect -300 -236 -292 -219
rect 292 -236 300 -219
rect 329 -236 337 -219
rect 921 -236 929 -219
rect 958 -236 966 -219
rect 1550 -236 1558 -219
rect -1638 -270 -1621 -239
rect 1621 -270 1638 -239
rect -1638 -287 -1590 -270
rect 1590 -287 1638 -270
<< viali >>
rect -1550 219 -966 236
rect -921 219 -337 236
rect -292 219 292 236
rect 337 219 921 236
rect 966 219 1550 236
rect -1581 -194 -1564 194
rect -952 -194 -935 194
rect -323 -194 -306 194
rect 306 -194 323 194
rect 935 -194 952 194
rect 1564 -194 1581 194
rect -1550 -236 -966 -219
rect -921 -236 -337 -219
rect -292 -236 292 -219
rect 337 -236 921 -219
rect 966 -236 1550 -219
<< metal1 >>
rect -1556 236 -960 239
rect -1556 219 -1550 236
rect -966 219 -960 236
rect -1556 216 -960 219
rect -927 236 -331 239
rect -927 219 -921 236
rect -337 219 -331 236
rect -927 216 -331 219
rect -298 236 298 239
rect -298 219 -292 236
rect 292 219 298 236
rect -298 216 298 219
rect 331 236 927 239
rect 331 219 337 236
rect 921 219 927 236
rect 331 216 927 219
rect 960 236 1556 239
rect 960 219 966 236
rect 1550 219 1556 236
rect 960 216 1556 219
rect -1584 194 -1561 200
rect -1584 -194 -1581 194
rect -1564 -194 -1561 194
rect -1584 -200 -1561 -194
rect -955 194 -932 200
rect -955 -194 -952 194
rect -935 -194 -932 194
rect -955 -200 -932 -194
rect -326 194 -303 200
rect -326 -194 -323 194
rect -306 -194 -303 194
rect -326 -200 -303 -194
rect 303 194 326 200
rect 303 -194 306 194
rect 323 -194 326 194
rect 303 -200 326 -194
rect 932 194 955 200
rect 932 -194 935 194
rect 952 -194 955 194
rect 932 -200 955 -194
rect 1561 194 1584 200
rect 1561 -194 1564 194
rect 1581 -194 1584 194
rect 1561 -200 1584 -194
rect -1556 -219 -960 -216
rect -1556 -236 -1550 -219
rect -966 -236 -960 -219
rect -1556 -239 -960 -236
rect -927 -219 -331 -216
rect -927 -236 -921 -219
rect -337 -236 -331 -219
rect -927 -239 -331 -236
rect -298 -219 298 -216
rect -298 -236 -292 -219
rect 292 -236 298 -219
rect -298 -239 298 -236
rect 331 -219 927 -216
rect 331 -236 337 -219
rect 921 -236 927 -219
rect 331 -239 927 -236
rect 960 -219 1556 -216
rect 960 -236 966 -219
rect 1550 -236 1556 -219
rect 960 -239 1556 -236
<< properties >>
string FIXED_BBOX -1629 -278 1629 278
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 4 l 6 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
