magic
tech sky130A
timestamp 1647254192
<< pwell >>
rect -2022 -186 2022 186
<< mvpsubdiff >>
rect -2004 162 -1668 168
rect -2004 145 -1950 162
rect -1722 145 -1668 162
rect -2004 139 -1668 145
rect -2004 114 -1975 139
rect -2004 -114 -1998 114
rect -1981 -114 -1975 114
rect -1697 114 -1668 139
rect -2004 -139 -1975 -114
rect -1697 -114 -1691 114
rect -1674 -114 -1668 114
rect -1697 -139 -1668 -114
rect -2004 -145 -1668 -139
rect -2004 -162 -1950 -145
rect -1722 -162 -1668 -145
rect -2004 -168 -1668 -162
rect -1596 162 -1260 168
rect -1596 145 -1542 162
rect -1314 145 -1260 162
rect -1596 139 -1260 145
rect -1596 114 -1567 139
rect -1596 -114 -1590 114
rect -1573 -114 -1567 114
rect -1289 114 -1260 139
rect -1596 -139 -1567 -114
rect -1289 -114 -1283 114
rect -1266 -114 -1260 114
rect -1289 -139 -1260 -114
rect -1596 -145 -1260 -139
rect -1596 -162 -1542 -145
rect -1314 -162 -1260 -145
rect -1596 -168 -1260 -162
rect -1188 162 -852 168
rect -1188 145 -1134 162
rect -906 145 -852 162
rect -1188 139 -852 145
rect -1188 114 -1159 139
rect -1188 -114 -1182 114
rect -1165 -114 -1159 114
rect -881 114 -852 139
rect -1188 -139 -1159 -114
rect -881 -114 -875 114
rect -858 -114 -852 114
rect -881 -139 -852 -114
rect -1188 -145 -852 -139
rect -1188 -162 -1134 -145
rect -906 -162 -852 -145
rect -1188 -168 -852 -162
rect -780 162 -444 168
rect -780 145 -726 162
rect -498 145 -444 162
rect -780 139 -444 145
rect -780 114 -751 139
rect -780 -114 -774 114
rect -757 -114 -751 114
rect -473 114 -444 139
rect -780 -139 -751 -114
rect -473 -114 -467 114
rect -450 -114 -444 114
rect -473 -139 -444 -114
rect -780 -145 -444 -139
rect -780 -162 -726 -145
rect -498 -162 -444 -145
rect -780 -168 -444 -162
rect -372 162 -36 168
rect -372 145 -318 162
rect -90 145 -36 162
rect -372 139 -36 145
rect -372 114 -343 139
rect -372 -114 -366 114
rect -349 -114 -343 114
rect -65 114 -36 139
rect -372 -139 -343 -114
rect -65 -114 -59 114
rect -42 -114 -36 114
rect -65 -139 -36 -114
rect -372 -145 -36 -139
rect -372 -162 -318 -145
rect -90 -162 -36 -145
rect -372 -168 -36 -162
rect 36 162 372 168
rect 36 145 90 162
rect 318 145 372 162
rect 36 139 372 145
rect 36 114 65 139
rect 36 -114 42 114
rect 59 -114 65 114
rect 343 114 372 139
rect 36 -139 65 -114
rect 343 -114 349 114
rect 366 -114 372 114
rect 343 -139 372 -114
rect 36 -145 372 -139
rect 36 -162 90 -145
rect 318 -162 372 -145
rect 36 -168 372 -162
rect 444 162 780 168
rect 444 145 498 162
rect 726 145 780 162
rect 444 139 780 145
rect 444 114 473 139
rect 444 -114 450 114
rect 467 -114 473 114
rect 751 114 780 139
rect 444 -139 473 -114
rect 751 -114 757 114
rect 774 -114 780 114
rect 751 -139 780 -114
rect 444 -145 780 -139
rect 444 -162 498 -145
rect 726 -162 780 -145
rect 444 -168 780 -162
rect 852 162 1188 168
rect 852 145 906 162
rect 1134 145 1188 162
rect 852 139 1188 145
rect 852 114 881 139
rect 852 -114 858 114
rect 875 -114 881 114
rect 1159 114 1188 139
rect 852 -139 881 -114
rect 1159 -114 1165 114
rect 1182 -114 1188 114
rect 1159 -139 1188 -114
rect 852 -145 1188 -139
rect 852 -162 906 -145
rect 1134 -162 1188 -145
rect 852 -168 1188 -162
rect 1260 162 1596 168
rect 1260 145 1314 162
rect 1542 145 1596 162
rect 1260 139 1596 145
rect 1260 114 1289 139
rect 1260 -114 1266 114
rect 1283 -114 1289 114
rect 1567 114 1596 139
rect 1260 -139 1289 -114
rect 1567 -114 1573 114
rect 1590 -114 1596 114
rect 1567 -139 1596 -114
rect 1260 -145 1596 -139
rect 1260 -162 1314 -145
rect 1542 -162 1596 -145
rect 1260 -168 1596 -162
rect 1668 162 2004 168
rect 1668 145 1722 162
rect 1950 145 2004 162
rect 1668 139 2004 145
rect 1668 114 1697 139
rect 1668 -114 1674 114
rect 1691 -114 1697 114
rect 1975 114 2004 139
rect 1668 -139 1697 -114
rect 1975 -114 1981 114
rect 1998 -114 2004 114
rect 1975 -139 2004 -114
rect 1668 -145 2004 -139
rect 1668 -162 1722 -145
rect 1950 -162 2004 -145
rect 1668 -168 2004 -162
<< mvpsubdiffcont >>
rect -1950 145 -1722 162
rect -1998 -114 -1981 114
rect -1691 -114 -1674 114
rect -1950 -162 -1722 -145
rect -1542 145 -1314 162
rect -1590 -114 -1573 114
rect -1283 -114 -1266 114
rect -1542 -162 -1314 -145
rect -1134 145 -906 162
rect -1182 -114 -1165 114
rect -875 -114 -858 114
rect -1134 -162 -906 -145
rect -726 145 -498 162
rect -774 -114 -757 114
rect -467 -114 -450 114
rect -726 -162 -498 -145
rect -318 145 -90 162
rect -366 -114 -349 114
rect -59 -114 -42 114
rect -318 -162 -90 -145
rect 90 145 318 162
rect 42 -114 59 114
rect 349 -114 366 114
rect 90 -162 318 -145
rect 498 145 726 162
rect 450 -114 467 114
rect 757 -114 774 114
rect 498 -162 726 -145
rect 906 145 1134 162
rect 858 -114 875 114
rect 1165 -114 1182 114
rect 906 -162 1134 -145
rect 1314 145 1542 162
rect 1266 -114 1283 114
rect 1573 -114 1590 114
rect 1314 -162 1542 -145
rect 1722 145 1950 162
rect 1674 -114 1691 114
rect 1981 -114 1998 114
rect 1722 -162 1950 -145
<< mvndiode >>
rect -1936 94 -1736 100
rect -1936 -94 -1930 94
rect -1742 -94 -1736 94
rect -1936 -100 -1736 -94
rect -1528 94 -1328 100
rect -1528 -94 -1522 94
rect -1334 -94 -1328 94
rect -1528 -100 -1328 -94
rect -1120 94 -920 100
rect -1120 -94 -1114 94
rect -926 -94 -920 94
rect -1120 -100 -920 -94
rect -712 94 -512 100
rect -712 -94 -706 94
rect -518 -94 -512 94
rect -712 -100 -512 -94
rect -304 94 -104 100
rect -304 -94 -298 94
rect -110 -94 -104 94
rect -304 -100 -104 -94
rect 104 94 304 100
rect 104 -94 110 94
rect 298 -94 304 94
rect 104 -100 304 -94
rect 512 94 712 100
rect 512 -94 518 94
rect 706 -94 712 94
rect 512 -100 712 -94
rect 920 94 1120 100
rect 920 -94 926 94
rect 1114 -94 1120 94
rect 920 -100 1120 -94
rect 1328 94 1528 100
rect 1328 -94 1334 94
rect 1522 -94 1528 94
rect 1328 -100 1528 -94
rect 1736 94 1936 100
rect 1736 -94 1742 94
rect 1930 -94 1936 94
rect 1736 -100 1936 -94
<< mvndiodec >>
rect -1930 -94 -1742 94
rect -1522 -94 -1334 94
rect -1114 -94 -926 94
rect -706 -94 -518 94
rect -298 -94 -110 94
rect 110 -94 298 94
rect 518 -94 706 94
rect 926 -94 1114 94
rect 1334 -94 1522 94
rect 1742 -94 1930 94
<< locali >>
rect -1998 145 -1950 162
rect -1722 145 -1674 162
rect -1998 114 -1981 145
rect -1691 114 -1674 145
rect -1938 -94 -1930 94
rect -1742 -94 -1734 94
rect -1998 -145 -1981 -114
rect -1691 -145 -1674 -114
rect -1998 -162 -1950 -145
rect -1722 -162 -1674 -145
rect -1590 145 -1542 162
rect -1314 145 -1266 162
rect -1590 114 -1573 145
rect -1283 114 -1266 145
rect -1530 -94 -1522 94
rect -1334 -94 -1326 94
rect -1590 -145 -1573 -114
rect -1283 -145 -1266 -114
rect -1590 -162 -1542 -145
rect -1314 -162 -1266 -145
rect -1182 145 -1134 162
rect -906 145 -858 162
rect -1182 114 -1165 145
rect -875 114 -858 145
rect -1122 -94 -1114 94
rect -926 -94 -918 94
rect -1182 -145 -1165 -114
rect -875 -145 -858 -114
rect -1182 -162 -1134 -145
rect -906 -162 -858 -145
rect -774 145 -726 162
rect -498 145 -450 162
rect -774 114 -757 145
rect -467 114 -450 145
rect -714 -94 -706 94
rect -518 -94 -510 94
rect -774 -145 -757 -114
rect -467 -145 -450 -114
rect -774 -162 -726 -145
rect -498 -162 -450 -145
rect -366 145 -318 162
rect -90 145 -42 162
rect -366 114 -349 145
rect -59 114 -42 145
rect -306 -94 -298 94
rect -110 -94 -102 94
rect -366 -145 -349 -114
rect -59 -145 -42 -114
rect -366 -162 -318 -145
rect -90 -162 -42 -145
rect 42 145 90 162
rect 318 145 366 162
rect 42 114 59 145
rect 349 114 366 145
rect 102 -94 110 94
rect 298 -94 306 94
rect 42 -145 59 -114
rect 349 -145 366 -114
rect 42 -162 90 -145
rect 318 -162 366 -145
rect 450 145 498 162
rect 726 145 774 162
rect 450 114 467 145
rect 757 114 774 145
rect 510 -94 518 94
rect 706 -94 714 94
rect 450 -145 467 -114
rect 757 -145 774 -114
rect 450 -162 498 -145
rect 726 -162 774 -145
rect 858 145 906 162
rect 1134 145 1182 162
rect 858 114 875 145
rect 1165 114 1182 145
rect 918 -94 926 94
rect 1114 -94 1122 94
rect 858 -145 875 -114
rect 1165 -145 1182 -114
rect 858 -162 906 -145
rect 1134 -162 1182 -145
rect 1266 145 1314 162
rect 1542 145 1590 162
rect 1266 114 1283 145
rect 1573 114 1590 145
rect 1326 -94 1334 94
rect 1522 -94 1530 94
rect 1266 -145 1283 -114
rect 1573 -145 1590 -114
rect 1266 -162 1314 -145
rect 1542 -162 1590 -145
rect 1674 145 1722 162
rect 1950 145 1998 162
rect 1674 114 1691 145
rect 1981 114 1998 145
rect 1734 -94 1742 94
rect 1930 -94 1938 94
rect 1674 -145 1691 -114
rect 1981 -145 1998 -114
rect 1674 -162 1722 -145
rect 1950 -162 1998 -145
<< viali >>
rect -1930 -94 -1742 94
rect -1522 -94 -1334 94
rect -1114 -94 -926 94
rect -706 -94 -518 94
rect -298 -94 -110 94
rect 110 -94 298 94
rect 518 -94 706 94
rect 926 -94 1114 94
rect 1334 -94 1522 94
rect 1742 -94 1930 94
<< metal1 >>
rect -1936 94 -1736 97
rect -1936 -94 -1930 94
rect -1742 -94 -1736 94
rect -1936 -97 -1736 -94
rect -1528 94 -1328 97
rect -1528 -94 -1522 94
rect -1334 -94 -1328 94
rect -1528 -97 -1328 -94
rect -1120 94 -920 97
rect -1120 -94 -1114 94
rect -926 -94 -920 94
rect -1120 -97 -920 -94
rect -712 94 -512 97
rect -712 -94 -706 94
rect -518 -94 -512 94
rect -712 -97 -512 -94
rect -304 94 -104 97
rect -304 -94 -298 94
rect -110 -94 -104 94
rect -304 -97 -104 -94
rect 104 94 304 97
rect 104 -94 110 94
rect 298 -94 304 94
rect 104 -97 304 -94
rect 512 94 712 97
rect 512 -94 518 94
rect 706 -94 712 94
rect 512 -97 712 -94
rect 920 94 1120 97
rect 920 -94 926 94
rect 1114 -94 1120 94
rect 920 -97 1120 -94
rect 1328 94 1528 97
rect 1328 -94 1334 94
rect 1522 -94 1528 94
rect 1328 -97 1528 -94
rect 1736 94 1936 97
rect 1736 -94 1742 94
rect 1930 -94 1936 94
rect 1736 -97 1936 -94
<< properties >>
string FIXED_BBOX 1682 -153 1989 153
string gencell sky130_fd_pr__diode_pw2nd_11v0
string library sky130
string parameters w 2 l 2 area 4.0 peri 8.0 nx 10 ny 1 dummy 0 lmin 0.45 wmin 0.45 elc 1 erc 1 etc 1 ebc 1 doverlap 0 compatible {sky130_fd_pr__diode_pw2nd_05v5 sky130_fd_pr__diode_pw2nd_05v5_lvt  sky130_fd_pr__diode_pw2nd_05v5_nvt sky130_fd_pr__diode_pw2nd_11v0} full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
