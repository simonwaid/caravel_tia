magic
tech sky130A
magscale 1 2
timestamp 1645787783
<< error_p >>
rect -715 599 -657 605
rect -519 599 -461 605
rect -323 599 -265 605
rect -127 599 -69 605
rect 69 599 127 605
rect 265 599 323 605
rect 461 599 519 605
rect 657 599 715 605
rect -715 565 -703 599
rect -519 565 -507 599
rect -323 565 -311 599
rect -127 565 -115 599
rect 69 565 81 599
rect 265 565 277 599
rect 461 565 473 599
rect 657 565 669 599
rect -715 559 -657 565
rect -519 559 -461 565
rect -323 559 -265 565
rect -127 559 -69 565
rect 69 559 127 565
rect 265 559 323 565
rect 461 559 519 565
rect 657 559 715 565
rect -617 71 -559 77
rect -421 71 -363 77
rect -225 71 -167 77
rect -29 71 29 77
rect 167 71 225 77
rect 363 71 421 77
rect 559 71 617 77
rect -617 37 -605 71
rect -421 37 -409 71
rect -225 37 -213 71
rect -29 37 -17 71
rect 167 37 179 71
rect 363 37 375 71
rect 559 37 571 71
rect -617 31 -559 37
rect -421 31 -363 37
rect -225 31 -167 37
rect -29 31 29 37
rect 167 31 225 37
rect 363 31 421 37
rect 559 31 617 37
rect -617 -37 -559 -31
rect -421 -37 -363 -31
rect -225 -37 -167 -31
rect -29 -37 29 -31
rect 167 -37 225 -31
rect 363 -37 421 -31
rect 559 -37 617 -31
rect -617 -71 -605 -37
rect -421 -71 -409 -37
rect -225 -71 -213 -37
rect -29 -71 -17 -37
rect 167 -71 179 -37
rect 363 -71 375 -37
rect 559 -71 571 -37
rect -617 -77 -559 -71
rect -421 -77 -363 -71
rect -225 -77 -167 -71
rect -29 -77 29 -71
rect 167 -77 225 -71
rect 363 -77 421 -71
rect 559 -77 617 -71
rect -715 -565 -657 -559
rect -519 -565 -461 -559
rect -323 -565 -265 -559
rect -127 -565 -69 -559
rect 69 -565 127 -559
rect 265 -565 323 -559
rect 461 -565 519 -559
rect 657 -565 715 -559
rect -715 -599 -703 -565
rect -519 -599 -507 -565
rect -323 -599 -311 -565
rect -127 -599 -115 -565
rect 69 -599 81 -565
rect 265 -599 277 -565
rect 461 -599 473 -565
rect 657 -599 669 -565
rect -715 -605 -657 -599
rect -519 -605 -461 -599
rect -323 -605 -265 -599
rect -127 -605 -69 -599
rect 69 -605 127 -599
rect 265 -605 323 -599
rect 461 -605 519 -599
rect 657 -605 715 -599
<< nwell >>
rect -902 -737 902 737
<< pmos >>
rect -706 118 -666 518
rect -608 118 -568 518
rect -510 118 -470 518
rect -412 118 -372 518
rect -314 118 -274 518
rect -216 118 -176 518
rect -118 118 -78 518
rect -20 118 20 518
rect 78 118 118 518
rect 176 118 216 518
rect 274 118 314 518
rect 372 118 412 518
rect 470 118 510 518
rect 568 118 608 518
rect 666 118 706 518
rect -706 -518 -666 -118
rect -608 -518 -568 -118
rect -510 -518 -470 -118
rect -412 -518 -372 -118
rect -314 -518 -274 -118
rect -216 -518 -176 -118
rect -118 -518 -78 -118
rect -20 -518 20 -118
rect 78 -518 118 -118
rect 176 -518 216 -118
rect 274 -518 314 -118
rect 372 -518 412 -118
rect 470 -518 510 -118
rect 568 -518 608 -118
rect 666 -518 706 -118
<< pdiff >>
rect -764 506 -706 518
rect -764 130 -752 506
rect -718 130 -706 506
rect -764 118 -706 130
rect -666 506 -608 518
rect -666 130 -654 506
rect -620 130 -608 506
rect -666 118 -608 130
rect -568 506 -510 518
rect -568 130 -556 506
rect -522 130 -510 506
rect -568 118 -510 130
rect -470 506 -412 518
rect -470 130 -458 506
rect -424 130 -412 506
rect -470 118 -412 130
rect -372 506 -314 518
rect -372 130 -360 506
rect -326 130 -314 506
rect -372 118 -314 130
rect -274 506 -216 518
rect -274 130 -262 506
rect -228 130 -216 506
rect -274 118 -216 130
rect -176 506 -118 518
rect -176 130 -164 506
rect -130 130 -118 506
rect -176 118 -118 130
rect -78 506 -20 518
rect -78 130 -66 506
rect -32 130 -20 506
rect -78 118 -20 130
rect 20 506 78 518
rect 20 130 32 506
rect 66 130 78 506
rect 20 118 78 130
rect 118 506 176 518
rect 118 130 130 506
rect 164 130 176 506
rect 118 118 176 130
rect 216 506 274 518
rect 216 130 228 506
rect 262 130 274 506
rect 216 118 274 130
rect 314 506 372 518
rect 314 130 326 506
rect 360 130 372 506
rect 314 118 372 130
rect 412 506 470 518
rect 412 130 424 506
rect 458 130 470 506
rect 412 118 470 130
rect 510 506 568 518
rect 510 130 522 506
rect 556 130 568 506
rect 510 118 568 130
rect 608 506 666 518
rect 608 130 620 506
rect 654 130 666 506
rect 608 118 666 130
rect 706 506 764 518
rect 706 130 718 506
rect 752 130 764 506
rect 706 118 764 130
rect -764 -130 -706 -118
rect -764 -506 -752 -130
rect -718 -506 -706 -130
rect -764 -518 -706 -506
rect -666 -130 -608 -118
rect -666 -506 -654 -130
rect -620 -506 -608 -130
rect -666 -518 -608 -506
rect -568 -130 -510 -118
rect -568 -506 -556 -130
rect -522 -506 -510 -130
rect -568 -518 -510 -506
rect -470 -130 -412 -118
rect -470 -506 -458 -130
rect -424 -506 -412 -130
rect -470 -518 -412 -506
rect -372 -130 -314 -118
rect -372 -506 -360 -130
rect -326 -506 -314 -130
rect -372 -518 -314 -506
rect -274 -130 -216 -118
rect -274 -506 -262 -130
rect -228 -506 -216 -130
rect -274 -518 -216 -506
rect -176 -130 -118 -118
rect -176 -506 -164 -130
rect -130 -506 -118 -130
rect -176 -518 -118 -506
rect -78 -130 -20 -118
rect -78 -506 -66 -130
rect -32 -506 -20 -130
rect -78 -518 -20 -506
rect 20 -130 78 -118
rect 20 -506 32 -130
rect 66 -506 78 -130
rect 20 -518 78 -506
rect 118 -130 176 -118
rect 118 -506 130 -130
rect 164 -506 176 -130
rect 118 -518 176 -506
rect 216 -130 274 -118
rect 216 -506 228 -130
rect 262 -506 274 -130
rect 216 -518 274 -506
rect 314 -130 372 -118
rect 314 -506 326 -130
rect 360 -506 372 -130
rect 314 -518 372 -506
rect 412 -130 470 -118
rect 412 -506 424 -130
rect 458 -506 470 -130
rect 412 -518 470 -506
rect 510 -130 568 -118
rect 510 -506 522 -130
rect 556 -506 568 -130
rect 510 -518 568 -506
rect 608 -130 666 -118
rect 608 -506 620 -130
rect 654 -506 666 -130
rect 608 -518 666 -506
rect 706 -130 764 -118
rect 706 -506 718 -130
rect 752 -506 764 -130
rect 706 -518 764 -506
<< pdiffc >>
rect -752 130 -718 506
rect -654 130 -620 506
rect -556 130 -522 506
rect -458 130 -424 506
rect -360 130 -326 506
rect -262 130 -228 506
rect -164 130 -130 506
rect -66 130 -32 506
rect 32 130 66 506
rect 130 130 164 506
rect 228 130 262 506
rect 326 130 360 506
rect 424 130 458 506
rect 522 130 556 506
rect 620 130 654 506
rect 718 130 752 506
rect -752 -506 -718 -130
rect -654 -506 -620 -130
rect -556 -506 -522 -130
rect -458 -506 -424 -130
rect -360 -506 -326 -130
rect -262 -506 -228 -130
rect -164 -506 -130 -130
rect -66 -506 -32 -130
rect 32 -506 66 -130
rect 130 -506 164 -130
rect 228 -506 262 -130
rect 326 -506 360 -130
rect 424 -506 458 -130
rect 522 -506 556 -130
rect 620 -506 654 -130
rect 718 -506 752 -130
<< nsubdiff >>
rect -866 667 -770 701
rect 770 667 866 701
rect -866 605 -832 667
rect 832 605 866 667
rect -866 -667 -832 -605
rect 832 -667 866 -605
rect -866 -701 -770 -667
rect 770 -701 866 -667
<< nsubdiffcont >>
rect -770 667 770 701
rect -866 -605 -832 605
rect 832 -605 866 605
rect -770 -701 770 -667
<< poly >>
rect -719 599 -653 615
rect -719 565 -703 599
rect -669 565 -653 599
rect -719 549 -653 565
rect -523 599 -457 615
rect -523 565 -507 599
rect -473 565 -457 599
rect -523 549 -457 565
rect -327 599 -261 615
rect -327 565 -311 599
rect -277 565 -261 599
rect -327 549 -261 565
rect -131 599 -65 615
rect -131 565 -115 599
rect -81 565 -65 599
rect -131 549 -65 565
rect 65 599 131 615
rect 65 565 81 599
rect 115 565 131 599
rect 65 549 131 565
rect 261 599 327 615
rect 261 565 277 599
rect 311 565 327 599
rect 261 549 327 565
rect 457 599 523 615
rect 457 565 473 599
rect 507 565 523 599
rect 457 549 523 565
rect 653 599 719 615
rect 653 565 669 599
rect 703 565 719 599
rect 653 549 719 565
rect -706 518 -666 549
rect -608 518 -568 544
rect -510 518 -470 549
rect -412 518 -372 544
rect -314 518 -274 549
rect -216 518 -176 544
rect -118 518 -78 549
rect -20 518 20 544
rect 78 518 118 549
rect 176 518 216 544
rect 274 518 314 549
rect 372 518 412 544
rect 470 518 510 549
rect 568 518 608 544
rect 666 518 706 549
rect -706 92 -666 118
rect -608 87 -568 118
rect -510 92 -470 118
rect -412 87 -372 118
rect -314 92 -274 118
rect -216 87 -176 118
rect -118 92 -78 118
rect -20 87 20 118
rect 78 92 118 118
rect 176 87 216 118
rect 274 92 314 118
rect 372 87 412 118
rect 470 92 510 118
rect 568 87 608 118
rect 666 92 706 118
rect -621 71 -555 87
rect -621 37 -605 71
rect -571 37 -555 71
rect -621 21 -555 37
rect -425 71 -359 87
rect -425 37 -409 71
rect -375 37 -359 71
rect -425 21 -359 37
rect -229 71 -163 87
rect -229 37 -213 71
rect -179 37 -163 71
rect -229 21 -163 37
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect 163 71 229 87
rect 163 37 179 71
rect 213 37 229 71
rect 163 21 229 37
rect 359 71 425 87
rect 359 37 375 71
rect 409 37 425 71
rect 359 21 425 37
rect 555 71 621 87
rect 555 37 571 71
rect 605 37 621 71
rect 555 21 621 37
rect -621 -37 -555 -21
rect -621 -71 -605 -37
rect -571 -71 -555 -37
rect -621 -87 -555 -71
rect -425 -37 -359 -21
rect -425 -71 -409 -37
rect -375 -71 -359 -37
rect -425 -87 -359 -71
rect -229 -37 -163 -21
rect -229 -71 -213 -37
rect -179 -71 -163 -37
rect -229 -87 -163 -71
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect 163 -37 229 -21
rect 163 -71 179 -37
rect 213 -71 229 -37
rect 163 -87 229 -71
rect 359 -37 425 -21
rect 359 -71 375 -37
rect 409 -71 425 -37
rect 359 -87 425 -71
rect 555 -37 621 -21
rect 555 -71 571 -37
rect 605 -71 621 -37
rect 555 -87 621 -71
rect -706 -118 -666 -92
rect -608 -118 -568 -87
rect -510 -118 -470 -92
rect -412 -118 -372 -87
rect -314 -118 -274 -92
rect -216 -118 -176 -87
rect -118 -118 -78 -92
rect -20 -118 20 -87
rect 78 -118 118 -92
rect 176 -118 216 -87
rect 274 -118 314 -92
rect 372 -118 412 -87
rect 470 -118 510 -92
rect 568 -118 608 -87
rect 666 -118 706 -92
rect -706 -549 -666 -518
rect -608 -544 -568 -518
rect -510 -549 -470 -518
rect -412 -544 -372 -518
rect -314 -549 -274 -518
rect -216 -544 -176 -518
rect -118 -549 -78 -518
rect -20 -544 20 -518
rect 78 -549 118 -518
rect 176 -544 216 -518
rect 274 -549 314 -518
rect 372 -544 412 -518
rect 470 -549 510 -518
rect 568 -544 608 -518
rect 666 -549 706 -518
rect -719 -565 -653 -549
rect -719 -599 -703 -565
rect -669 -599 -653 -565
rect -719 -615 -653 -599
rect -523 -565 -457 -549
rect -523 -599 -507 -565
rect -473 -599 -457 -565
rect -523 -615 -457 -599
rect -327 -565 -261 -549
rect -327 -599 -311 -565
rect -277 -599 -261 -565
rect -327 -615 -261 -599
rect -131 -565 -65 -549
rect -131 -599 -115 -565
rect -81 -599 -65 -565
rect -131 -615 -65 -599
rect 65 -565 131 -549
rect 65 -599 81 -565
rect 115 -599 131 -565
rect 65 -615 131 -599
rect 261 -565 327 -549
rect 261 -599 277 -565
rect 311 -599 327 -565
rect 261 -615 327 -599
rect 457 -565 523 -549
rect 457 -599 473 -565
rect 507 -599 523 -565
rect 457 -615 523 -599
rect 653 -565 719 -549
rect 653 -599 669 -565
rect 703 -599 719 -565
rect 653 -615 719 -599
<< polycont >>
rect -703 565 -669 599
rect -507 565 -473 599
rect -311 565 -277 599
rect -115 565 -81 599
rect 81 565 115 599
rect 277 565 311 599
rect 473 565 507 599
rect 669 565 703 599
rect -605 37 -571 71
rect -409 37 -375 71
rect -213 37 -179 71
rect -17 37 17 71
rect 179 37 213 71
rect 375 37 409 71
rect 571 37 605 71
rect -605 -71 -571 -37
rect -409 -71 -375 -37
rect -213 -71 -179 -37
rect -17 -71 17 -37
rect 179 -71 213 -37
rect 375 -71 409 -37
rect 571 -71 605 -37
rect -703 -599 -669 -565
rect -507 -599 -473 -565
rect -311 -599 -277 -565
rect -115 -599 -81 -565
rect 81 -599 115 -565
rect 277 -599 311 -565
rect 473 -599 507 -565
rect 669 -599 703 -565
<< locali >>
rect -866 667 -770 701
rect 770 667 866 701
rect -866 605 -832 667
rect 832 605 866 667
rect -719 565 -703 599
rect -669 565 -653 599
rect -523 565 -507 599
rect -473 565 -457 599
rect -327 565 -311 599
rect -277 565 -261 599
rect -131 565 -115 599
rect -81 565 -65 599
rect 65 565 81 599
rect 115 565 131 599
rect 261 565 277 599
rect 311 565 327 599
rect 457 565 473 599
rect 507 565 523 599
rect 653 565 669 599
rect 703 565 719 599
rect -752 506 -718 522
rect -752 114 -718 130
rect -654 506 -620 522
rect -654 114 -620 130
rect -556 506 -522 522
rect -556 114 -522 130
rect -458 506 -424 522
rect -458 114 -424 130
rect -360 506 -326 522
rect -360 114 -326 130
rect -262 506 -228 522
rect -262 114 -228 130
rect -164 506 -130 522
rect -164 114 -130 130
rect -66 506 -32 522
rect -66 114 -32 130
rect 32 506 66 522
rect 32 114 66 130
rect 130 506 164 522
rect 130 114 164 130
rect 228 506 262 522
rect 228 114 262 130
rect 326 506 360 522
rect 326 114 360 130
rect 424 506 458 522
rect 424 114 458 130
rect 522 506 556 522
rect 522 114 556 130
rect 620 506 654 522
rect 620 114 654 130
rect 718 506 752 522
rect 718 114 752 130
rect -621 37 -605 71
rect -571 37 -555 71
rect -425 37 -409 71
rect -375 37 -359 71
rect -229 37 -213 71
rect -179 37 -163 71
rect -33 37 -17 71
rect 17 37 33 71
rect 163 37 179 71
rect 213 37 229 71
rect 359 37 375 71
rect 409 37 425 71
rect 555 37 571 71
rect 605 37 621 71
rect -621 -71 -605 -37
rect -571 -71 -555 -37
rect -425 -71 -409 -37
rect -375 -71 -359 -37
rect -229 -71 -213 -37
rect -179 -71 -163 -37
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect 163 -71 179 -37
rect 213 -71 229 -37
rect 359 -71 375 -37
rect 409 -71 425 -37
rect 555 -71 571 -37
rect 605 -71 621 -37
rect -752 -130 -718 -114
rect -752 -522 -718 -506
rect -654 -130 -620 -114
rect -654 -522 -620 -506
rect -556 -130 -522 -114
rect -556 -522 -522 -506
rect -458 -130 -424 -114
rect -458 -522 -424 -506
rect -360 -130 -326 -114
rect -360 -522 -326 -506
rect -262 -130 -228 -114
rect -262 -522 -228 -506
rect -164 -130 -130 -114
rect -164 -522 -130 -506
rect -66 -130 -32 -114
rect -66 -522 -32 -506
rect 32 -130 66 -114
rect 32 -522 66 -506
rect 130 -130 164 -114
rect 130 -522 164 -506
rect 228 -130 262 -114
rect 228 -522 262 -506
rect 326 -130 360 -114
rect 326 -522 360 -506
rect 424 -130 458 -114
rect 424 -522 458 -506
rect 522 -130 556 -114
rect 522 -522 556 -506
rect 620 -130 654 -114
rect 620 -522 654 -506
rect 718 -130 752 -114
rect 718 -522 752 -506
rect -719 -599 -703 -565
rect -669 -599 -653 -565
rect -523 -599 -507 -565
rect -473 -599 -457 -565
rect -327 -599 -311 -565
rect -277 -599 -261 -565
rect -131 -599 -115 -565
rect -81 -599 -65 -565
rect 65 -599 81 -565
rect 115 -599 131 -565
rect 261 -599 277 -565
rect 311 -599 327 -565
rect 457 -599 473 -565
rect 507 -599 523 -565
rect 653 -599 669 -565
rect 703 -599 719 -565
rect -866 -667 -832 -605
rect 832 -667 866 -605
rect -866 -701 -770 -667
rect 770 -701 866 -667
<< viali >>
rect -703 565 -669 599
rect -507 565 -473 599
rect -311 565 -277 599
rect -115 565 -81 599
rect 81 565 115 599
rect 277 565 311 599
rect 473 565 507 599
rect 669 565 703 599
rect -752 130 -718 506
rect -654 130 -620 506
rect -556 130 -522 506
rect -458 130 -424 506
rect -360 130 -326 506
rect -262 130 -228 506
rect -164 130 -130 506
rect -66 130 -32 506
rect 32 130 66 506
rect 130 130 164 506
rect 228 130 262 506
rect 326 130 360 506
rect 424 130 458 506
rect 522 130 556 506
rect 620 130 654 506
rect 718 130 752 506
rect -605 37 -571 71
rect -409 37 -375 71
rect -213 37 -179 71
rect -17 37 17 71
rect 179 37 213 71
rect 375 37 409 71
rect 571 37 605 71
rect -605 -71 -571 -37
rect -409 -71 -375 -37
rect -213 -71 -179 -37
rect -17 -71 17 -37
rect 179 -71 213 -37
rect 375 -71 409 -37
rect 571 -71 605 -37
rect -752 -506 -718 -130
rect -654 -506 -620 -130
rect -556 -506 -522 -130
rect -458 -506 -424 -130
rect -360 -506 -326 -130
rect -262 -506 -228 -130
rect -164 -506 -130 -130
rect -66 -506 -32 -130
rect 32 -506 66 -130
rect 130 -506 164 -130
rect 228 -506 262 -130
rect 326 -506 360 -130
rect 424 -506 458 -130
rect 522 -506 556 -130
rect 620 -506 654 -130
rect 718 -506 752 -130
rect -703 -599 -669 -565
rect -507 -599 -473 -565
rect -311 -599 -277 -565
rect -115 -599 -81 -565
rect 81 -599 115 -565
rect 277 -599 311 -565
rect 473 -599 507 -565
rect 669 -599 703 -565
<< metal1 >>
rect -715 599 -657 605
rect -715 565 -703 599
rect -669 565 -657 599
rect -715 559 -657 565
rect -519 599 -461 605
rect -519 565 -507 599
rect -473 565 -461 599
rect -519 559 -461 565
rect -323 599 -265 605
rect -323 565 -311 599
rect -277 565 -265 599
rect -323 559 -265 565
rect -127 599 -69 605
rect -127 565 -115 599
rect -81 565 -69 599
rect -127 559 -69 565
rect 69 599 127 605
rect 69 565 81 599
rect 115 565 127 599
rect 69 559 127 565
rect 265 599 323 605
rect 265 565 277 599
rect 311 565 323 599
rect 265 559 323 565
rect 461 599 519 605
rect 461 565 473 599
rect 507 565 519 599
rect 461 559 519 565
rect 657 599 715 605
rect 657 565 669 599
rect 703 565 715 599
rect 657 559 715 565
rect -758 506 -712 518
rect -758 130 -752 506
rect -718 130 -712 506
rect -758 118 -712 130
rect -660 506 -614 518
rect -660 130 -654 506
rect -620 130 -614 506
rect -660 118 -614 130
rect -562 506 -516 518
rect -562 130 -556 506
rect -522 130 -516 506
rect -562 118 -516 130
rect -464 506 -418 518
rect -464 130 -458 506
rect -424 130 -418 506
rect -464 118 -418 130
rect -366 506 -320 518
rect -366 130 -360 506
rect -326 130 -320 506
rect -366 118 -320 130
rect -268 506 -222 518
rect -268 130 -262 506
rect -228 130 -222 506
rect -268 118 -222 130
rect -170 506 -124 518
rect -170 130 -164 506
rect -130 130 -124 506
rect -170 118 -124 130
rect -72 506 -26 518
rect -72 130 -66 506
rect -32 130 -26 506
rect -72 118 -26 130
rect 26 506 72 518
rect 26 130 32 506
rect 66 130 72 506
rect 26 118 72 130
rect 124 506 170 518
rect 124 130 130 506
rect 164 130 170 506
rect 124 118 170 130
rect 222 506 268 518
rect 222 130 228 506
rect 262 130 268 506
rect 222 118 268 130
rect 320 506 366 518
rect 320 130 326 506
rect 360 130 366 506
rect 320 118 366 130
rect 418 506 464 518
rect 418 130 424 506
rect 458 130 464 506
rect 418 118 464 130
rect 516 506 562 518
rect 516 130 522 506
rect 556 130 562 506
rect 516 118 562 130
rect 614 506 660 518
rect 614 130 620 506
rect 654 130 660 506
rect 614 118 660 130
rect 712 506 758 518
rect 712 130 718 506
rect 752 130 758 506
rect 712 118 758 130
rect -617 71 -559 77
rect -617 37 -605 71
rect -571 37 -559 71
rect -617 31 -559 37
rect -421 71 -363 77
rect -421 37 -409 71
rect -375 37 -363 71
rect -421 31 -363 37
rect -225 71 -167 77
rect -225 37 -213 71
rect -179 37 -167 71
rect -225 31 -167 37
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect 167 71 225 77
rect 167 37 179 71
rect 213 37 225 71
rect 167 31 225 37
rect 363 71 421 77
rect 363 37 375 71
rect 409 37 421 71
rect 363 31 421 37
rect 559 71 617 77
rect 559 37 571 71
rect 605 37 617 71
rect 559 31 617 37
rect -617 -37 -559 -31
rect -617 -71 -605 -37
rect -571 -71 -559 -37
rect -617 -77 -559 -71
rect -421 -37 -363 -31
rect -421 -71 -409 -37
rect -375 -71 -363 -37
rect -421 -77 -363 -71
rect -225 -37 -167 -31
rect -225 -71 -213 -37
rect -179 -71 -167 -37
rect -225 -77 -167 -71
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect 167 -37 225 -31
rect 167 -71 179 -37
rect 213 -71 225 -37
rect 167 -77 225 -71
rect 363 -37 421 -31
rect 363 -71 375 -37
rect 409 -71 421 -37
rect 363 -77 421 -71
rect 559 -37 617 -31
rect 559 -71 571 -37
rect 605 -71 617 -37
rect 559 -77 617 -71
rect -758 -130 -712 -118
rect -758 -506 -752 -130
rect -718 -506 -712 -130
rect -758 -518 -712 -506
rect -660 -130 -614 -118
rect -660 -506 -654 -130
rect -620 -506 -614 -130
rect -660 -518 -614 -506
rect -562 -130 -516 -118
rect -562 -506 -556 -130
rect -522 -506 -516 -130
rect -562 -518 -516 -506
rect -464 -130 -418 -118
rect -464 -506 -458 -130
rect -424 -506 -418 -130
rect -464 -518 -418 -506
rect -366 -130 -320 -118
rect -366 -506 -360 -130
rect -326 -506 -320 -130
rect -366 -518 -320 -506
rect -268 -130 -222 -118
rect -268 -506 -262 -130
rect -228 -506 -222 -130
rect -268 -518 -222 -506
rect -170 -130 -124 -118
rect -170 -506 -164 -130
rect -130 -506 -124 -130
rect -170 -518 -124 -506
rect -72 -130 -26 -118
rect -72 -506 -66 -130
rect -32 -506 -26 -130
rect -72 -518 -26 -506
rect 26 -130 72 -118
rect 26 -506 32 -130
rect 66 -506 72 -130
rect 26 -518 72 -506
rect 124 -130 170 -118
rect 124 -506 130 -130
rect 164 -506 170 -130
rect 124 -518 170 -506
rect 222 -130 268 -118
rect 222 -506 228 -130
rect 262 -506 268 -130
rect 222 -518 268 -506
rect 320 -130 366 -118
rect 320 -506 326 -130
rect 360 -506 366 -130
rect 320 -518 366 -506
rect 418 -130 464 -118
rect 418 -506 424 -130
rect 458 -506 464 -130
rect 418 -518 464 -506
rect 516 -130 562 -118
rect 516 -506 522 -130
rect 556 -506 562 -130
rect 516 -518 562 -506
rect 614 -130 660 -118
rect 614 -506 620 -130
rect 654 -506 660 -130
rect 614 -518 660 -506
rect 712 -130 758 -118
rect 712 -506 718 -130
rect 752 -506 758 -130
rect 712 -518 758 -506
rect -715 -565 -657 -559
rect -715 -599 -703 -565
rect -669 -599 -657 -565
rect -715 -605 -657 -599
rect -519 -565 -461 -559
rect -519 -599 -507 -565
rect -473 -599 -461 -565
rect -519 -605 -461 -599
rect -323 -565 -265 -559
rect -323 -599 -311 -565
rect -277 -599 -265 -565
rect -323 -605 -265 -599
rect -127 -565 -69 -559
rect -127 -599 -115 -565
rect -81 -599 -69 -565
rect -127 -605 -69 -599
rect 69 -565 127 -559
rect 69 -599 81 -565
rect 115 -599 127 -565
rect 69 -605 127 -599
rect 265 -565 323 -559
rect 265 -599 277 -565
rect 311 -599 323 -565
rect 265 -605 323 -599
rect 461 -565 519 -559
rect 461 -599 473 -565
rect 507 -599 519 -565
rect 461 -605 519 -599
rect 657 -565 715 -559
rect 657 -599 669 -565
rect 703 -599 715 -565
rect 657 -605 715 -599
<< properties >>
string FIXED_BBOX -849 -684 849 684
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 0.2 m 2 nf 15 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
