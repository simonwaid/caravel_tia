magic
tech sky130A
magscale 1 2
timestamp 1646401284
<< nwell >>
rect 230 1520 310 1570
<< locali >>
rect -320 1630 410 1700
rect -320 910 -260 1630
rect 340 910 410 1630
rect -320 870 410 910
rect -320 820 1050 870
rect -320 -1820 -160 820
rect 340 810 1050 820
rect 890 -1820 1050 810
rect -320 -1880 1050 -1820
<< metal1 >>
rect -40 1520 390 1590
rect -190 1320 -180 1480
rect -126 1320 -116 1480
rect 6 1320 16 1480
rect 70 1320 80 1480
rect 202 1320 212 1480
rect 266 1320 276 1480
rect -92 1078 -82 1238
rect -28 1078 -18 1238
rect 104 1078 114 1238
rect 168 1078 178 1238
rect 310 1040 390 1520
rect -140 970 390 1040
rect -70 740 10 970
rect -130 690 860 740
rect -190 488 -180 648
rect -126 488 -116 648
rect -70 210 10 690
rect 326 488 336 648
rect 390 488 400 648
rect 842 488 852 648
rect 906 488 916 648
rect 68 246 78 406
rect 132 246 142 406
rect 584 246 594 406
rect 648 246 658 406
rect -130 50 860 210
rect -190 -390 -180 -230
rect -126 -390 -116 -230
rect -70 -430 10 50
rect 68 -148 78 12
rect 132 -148 142 12
rect 584 -148 594 12
rect 648 -148 658 12
rect 326 -390 336 -230
rect 390 -390 400 -230
rect 842 -390 852 -230
rect 906 -390 916 -230
rect -130 -590 860 -430
rect -190 -784 -180 -624
rect -126 -784 -116 -624
rect -70 -1060 10 -590
rect 326 -784 336 -624
rect 390 -784 400 -624
rect 842 -784 852 -624
rect 906 -784 916 -624
rect 68 -1026 78 -866
rect 132 -1026 142 -866
rect 584 -1026 594 -866
rect 648 -1026 658 -866
rect -130 -1220 860 -1060
rect -190 -1662 -180 -1502
rect -126 -1662 -116 -1502
rect -70 -1700 10 -1220
rect 68 -1420 78 -1260
rect 132 -1420 142 -1260
rect 584 -1420 594 -1260
rect 648 -1420 658 -1260
rect 326 -1662 336 -1502
rect 390 -1662 400 -1502
rect 842 -1662 852 -1502
rect 906 -1662 916 -1502
rect -130 -1750 860 -1700
<< via1 >>
rect -180 1320 -126 1480
rect 16 1320 70 1480
rect 212 1320 266 1480
rect -82 1078 -28 1238
rect 114 1078 168 1238
rect -180 488 -126 648
rect 336 488 390 648
rect 852 488 906 648
rect 78 246 132 406
rect 594 246 648 406
rect -180 -390 -126 -230
rect 78 -148 132 12
rect 594 -148 648 12
rect 336 -390 390 -230
rect 852 -390 906 -230
rect -180 -784 -126 -624
rect 336 -784 390 -624
rect 852 -784 906 -624
rect 78 -1026 132 -866
rect 594 -1026 648 -866
rect -180 -1662 -126 -1502
rect 78 -1420 132 -1260
rect 594 -1420 648 -1260
rect 336 -1662 390 -1502
rect 852 -1662 906 -1502
<< metal2 >>
rect -190 1480 270 1490
rect -190 1320 -180 1480
rect -126 1320 16 1480
rect 70 1320 212 1480
rect 266 1320 270 1480
rect -190 1300 270 1320
rect 70 1250 650 1260
rect -90 1238 70 1250
rect -90 1078 -82 1238
rect -28 1078 70 1238
rect -90 1060 70 1078
rect 70 1050 650 1060
rect -240 650 960 660
rect 0 648 720 650
rect 0 488 336 648
rect 390 488 720 648
rect 0 480 720 488
rect -240 470 960 480
rect 70 410 650 420
rect 70 406 80 410
rect 640 406 650 410
rect 70 246 78 406
rect 648 246 650 406
rect 70 240 80 246
rect 640 240 650 246
rect 70 230 650 240
rect 70 20 650 30
rect 70 12 80 20
rect 640 12 650 20
rect 70 -148 78 12
rect 648 -148 650 12
rect 70 -150 80 -148
rect 640 -150 650 -148
rect 70 -160 650 -150
rect -240 -230 960 -220
rect 0 -390 336 -230
rect 390 -390 720 -230
rect 0 -400 720 -390
rect -240 -410 960 -400
rect -240 -620 960 -610
rect 0 -624 720 -620
rect 0 -784 336 -624
rect 390 -784 720 -624
rect 0 -790 720 -784
rect -240 -800 960 -790
rect 70 -860 660 -850
rect 70 -866 80 -860
rect 640 -866 660 -860
rect 70 -1026 78 -866
rect 648 -1026 660 -866
rect 70 -1030 80 -1026
rect 640 -1030 660 -1026
rect 70 -1040 660 -1030
rect 70 -1260 650 -1250
rect 70 -1420 78 -1260
rect 648 -1420 650 -1260
rect 70 -1430 80 -1420
rect 640 -1430 650 -1420
rect 70 -1440 650 -1430
rect -240 -1500 960 -1490
rect 0 -1502 720 -1500
rect 0 -1662 336 -1502
rect 390 -1662 720 -1502
rect 0 -1670 720 -1662
rect -240 -1680 960 -1670
<< via2 >>
rect 70 1238 650 1250
rect 70 1078 114 1238
rect 114 1078 168 1238
rect 168 1078 650 1238
rect 70 1060 650 1078
rect -240 648 0 650
rect 720 648 960 650
rect -240 488 -180 648
rect -180 488 -126 648
rect -126 488 0 648
rect 720 488 852 648
rect 852 488 906 648
rect 906 488 960 648
rect -240 480 0 488
rect 720 480 960 488
rect 80 406 640 410
rect 80 246 132 406
rect 132 246 594 406
rect 594 246 640 406
rect 80 240 640 246
rect 80 12 640 20
rect 80 -148 132 12
rect 132 -148 594 12
rect 594 -148 640 12
rect 80 -150 640 -148
rect -240 -390 -180 -230
rect -180 -390 -126 -230
rect -126 -390 0 -230
rect 720 -390 852 -230
rect 852 -390 906 -230
rect 906 -390 960 -230
rect -240 -400 0 -390
rect 720 -400 960 -390
rect -240 -624 0 -620
rect 720 -624 960 -620
rect -240 -784 -180 -624
rect -180 -784 -126 -624
rect -126 -784 0 -624
rect 720 -784 852 -624
rect 852 -784 906 -624
rect 906 -784 960 -624
rect -240 -790 0 -784
rect 720 -790 960 -784
rect 80 -866 640 -860
rect 80 -1026 132 -866
rect 132 -1026 594 -866
rect 594 -1026 640 -866
rect 80 -1030 640 -1026
rect 80 -1420 132 -1260
rect 132 -1420 594 -1260
rect 594 -1420 640 -1260
rect 80 -1430 640 -1420
rect -240 -1502 0 -1500
rect 720 -1502 960 -1500
rect -240 -1662 -180 -1502
rect -180 -1662 -126 -1502
rect -126 -1662 0 -1502
rect 720 -1662 852 -1502
rect 852 -1662 906 -1502
rect 906 -1662 960 -1502
rect -240 -1670 0 -1662
rect 720 -1670 960 -1662
<< metal3 >>
rect 60 1250 660 1255
rect 60 1060 70 1250
rect 650 1060 660 1250
rect 60 1055 660 1060
rect -230 655 10 660
rect -250 650 10 655
rect -250 480 -240 650
rect 0 480 10 650
rect -250 475 10 480
rect -230 -225 10 475
rect -250 -230 10 -225
rect -250 -400 -240 -230
rect 0 -400 10 -230
rect -250 -405 10 -400
rect -230 -615 10 -405
rect -250 -620 10 -615
rect -250 -790 -240 -620
rect 0 -790 10 -620
rect -250 -795 10 -790
rect -230 -1495 10 -795
rect 70 410 650 1055
rect 70 240 80 410
rect 640 240 650 410
rect 70 20 650 240
rect 70 -150 80 20
rect 640 -150 650 20
rect 70 -860 650 -150
rect 70 -1030 80 -860
rect 640 -1030 650 -860
rect 70 -1260 650 -1030
rect 70 -1430 80 -1260
rect 640 -1430 650 -1260
rect 70 -1440 650 -1430
rect 710 655 960 660
rect 710 650 970 655
rect 710 480 720 650
rect 960 480 970 650
rect 710 475 970 480
rect 710 -225 960 475
rect 710 -230 970 -225
rect 710 -400 720 -230
rect 960 -400 970 -230
rect 710 -405 970 -400
rect 710 -615 960 -405
rect 710 -620 970 -615
rect 710 -790 720 -620
rect 960 -790 970 -620
rect 710 -795 970 -790
rect -250 -1500 10 -1495
rect -250 -1670 -240 -1500
rect 0 -1540 10 -1500
rect 710 -1495 960 -795
rect 710 -1500 970 -1495
rect 710 -1540 720 -1500
rect 0 -1670 720 -1540
rect 960 -1670 970 -1500
rect -250 -1675 970 -1670
rect -230 -1880 960 -1675
use sky130_fd_pr__pfet_01v8_LXX5YL  sky130_fd_pr__pfet_01v8_LXX5YL_0
timestamp 1646400034
transform 1 0 363 0 1 -507
box -683 -1373 683 1373
use sky130_fd_pr__pfet_01v8_X9CJL2  sky130_fd_pr__pfet_01v8_X9CJL2_0
timestamp 1646401284
transform 1 0 43 0 1 1279
box -363 -419 363 419
<< end >>
