magic
tech sky130A
magscale 1 2
timestamp 1646921651
<< pwell >>
rect 2 2306 1508 2372
rect 2 1796 1508 1862
rect 2 1688 1508 1754
rect 2 1178 1508 1244
rect 2 1070 1508 1136
rect 2 560 1508 626
rect 2 452 1508 518
rect 2 -58 1508 8
<< poly >>
rect 2 2356 1508 2372
rect 2 2322 114 2356
rect 148 2322 306 2356
rect 340 2322 498 2356
rect 532 2322 690 2356
rect 724 2322 882 2356
rect 916 2322 1074 2356
rect 1108 2322 1266 2356
rect 1300 2322 1458 2356
rect 1492 2322 1508 2356
rect 2 2306 1508 2322
rect 2 1846 1508 1862
rect 2 1812 18 1846
rect 52 1812 210 1846
rect 244 1812 402 1846
rect 436 1812 594 1846
rect 628 1812 786 1846
rect 820 1812 978 1846
rect 1012 1812 1170 1846
rect 1204 1812 1362 1846
rect 1396 1812 1508 1846
rect 2 1796 1508 1812
rect 2 1738 1508 1754
rect 2 1704 18 1738
rect 52 1704 210 1738
rect 244 1704 402 1738
rect 436 1704 594 1738
rect 628 1704 786 1738
rect 820 1704 978 1738
rect 1012 1704 1170 1738
rect 1204 1704 1362 1738
rect 1396 1704 1508 1738
rect 2 1688 1508 1704
rect 2 1228 1508 1244
rect 2 1194 114 1228
rect 148 1194 306 1228
rect 340 1194 498 1228
rect 532 1194 690 1228
rect 724 1194 882 1228
rect 916 1194 1074 1228
rect 1108 1194 1266 1228
rect 1300 1194 1458 1228
rect 1492 1194 1508 1228
rect 2 1178 1508 1194
rect 2 1120 1508 1136
rect 2 1086 114 1120
rect 148 1086 306 1120
rect 340 1086 498 1120
rect 532 1086 690 1120
rect 724 1086 882 1120
rect 916 1086 1074 1120
rect 1108 1086 1266 1120
rect 1300 1086 1458 1120
rect 1492 1086 1508 1120
rect 2 1070 1508 1086
rect 2 610 1508 626
rect 2 576 18 610
rect 52 576 210 610
rect 244 576 402 610
rect 436 576 594 610
rect 628 576 786 610
rect 820 576 978 610
rect 1012 576 1170 610
rect 1204 576 1362 610
rect 1396 576 1508 610
rect 2 560 1508 576
rect 2 502 1508 518
rect 2 468 18 502
rect 52 468 210 502
rect 244 468 402 502
rect 436 468 594 502
rect 628 468 786 502
rect 820 468 978 502
rect 1012 468 1170 502
rect 1204 468 1362 502
rect 1396 468 1508 502
rect 2 452 1508 468
rect 2 -8 1508 8
rect 2 -42 114 -8
rect 148 -42 306 -8
rect 340 -42 498 -8
rect 532 -42 690 -8
rect 724 -42 882 -8
rect 916 -42 1074 -8
rect 1108 -42 1266 -8
rect 1300 -42 1458 -8
rect 1492 -42 1508 -8
rect 2 -58 1508 -42
<< polycont >>
rect 114 2322 148 2356
rect 306 2322 340 2356
rect 498 2322 532 2356
rect 690 2322 724 2356
rect 882 2322 916 2356
rect 1074 2322 1108 2356
rect 1266 2322 1300 2356
rect 1458 2322 1492 2356
rect 18 1812 52 1846
rect 210 1812 244 1846
rect 402 1812 436 1846
rect 594 1812 628 1846
rect 786 1812 820 1846
rect 978 1812 1012 1846
rect 1170 1812 1204 1846
rect 1362 1812 1396 1846
rect 18 1704 52 1738
rect 210 1704 244 1738
rect 402 1704 436 1738
rect 594 1704 628 1738
rect 786 1704 820 1738
rect 978 1704 1012 1738
rect 1170 1704 1204 1738
rect 1362 1704 1396 1738
rect 114 1194 148 1228
rect 306 1194 340 1228
rect 498 1194 532 1228
rect 690 1194 724 1228
rect 882 1194 916 1228
rect 1074 1194 1108 1228
rect 1266 1194 1300 1228
rect 1458 1194 1492 1228
rect 114 1086 148 1120
rect 306 1086 340 1120
rect 498 1086 532 1120
rect 690 1086 724 1120
rect 882 1086 916 1120
rect 1074 1086 1108 1120
rect 1266 1086 1300 1120
rect 1458 1086 1492 1120
rect 18 576 52 610
rect 210 576 244 610
rect 402 576 436 610
rect 594 576 628 610
rect 786 576 820 610
rect 978 576 1012 610
rect 1170 576 1204 610
rect 1362 576 1396 610
rect 18 468 52 502
rect 210 468 244 502
rect 402 468 436 502
rect 594 468 628 502
rect 786 468 820 502
rect 978 468 1012 502
rect 1170 468 1204 502
rect 1362 468 1396 502
rect 114 -42 148 -8
rect 306 -42 340 -8
rect 498 -42 532 -8
rect 690 -42 724 -8
rect 882 -42 916 -8
rect 1074 -42 1108 -8
rect 1266 -42 1300 -8
rect 1458 -42 1492 -8
<< locali >>
rect 2 2322 114 2356
rect 148 2322 306 2356
rect 340 2322 498 2356
rect 532 2322 690 2356
rect 724 2322 882 2356
rect 916 2322 1074 2356
rect 1108 2322 1266 2356
rect 1300 2322 1458 2356
rect 1492 2322 1508 2356
rect 2 1812 18 1846
rect 52 1812 210 1846
rect 244 1812 402 1846
rect 436 1812 594 1846
rect 628 1812 786 1846
rect 820 1812 978 1846
rect 1012 1812 1170 1846
rect 1204 1812 1362 1846
rect 1396 1812 1508 1846
rect 2 1704 18 1738
rect 52 1704 210 1738
rect 244 1704 402 1738
rect 436 1704 594 1738
rect 628 1704 786 1738
rect 820 1704 978 1738
rect 1012 1704 1170 1738
rect 1204 1704 1362 1738
rect 1396 1704 1508 1738
rect 2 1194 114 1228
rect 148 1194 306 1228
rect 340 1194 498 1228
rect 532 1194 690 1228
rect 724 1194 882 1228
rect 916 1194 1074 1228
rect 1108 1194 1266 1228
rect 1300 1194 1458 1228
rect 1492 1194 1508 1228
rect 2 1086 114 1120
rect 148 1086 306 1120
rect 340 1086 498 1120
rect 532 1086 690 1120
rect 724 1086 882 1120
rect 916 1086 1074 1120
rect 1108 1086 1266 1120
rect 1300 1086 1458 1120
rect 1492 1086 1508 1120
rect 2 576 18 610
rect 52 576 210 610
rect 244 576 402 610
rect 436 576 594 610
rect 628 576 786 610
rect 820 576 978 610
rect 1012 576 1170 610
rect 1204 576 1362 610
rect 1396 576 1508 610
rect 2 468 18 502
rect 52 468 210 502
rect 244 468 402 502
rect 436 468 594 502
rect 628 468 786 502
rect 820 468 978 502
rect 1012 468 1170 502
rect 1204 468 1362 502
rect 1396 468 1508 502
rect 2 -42 114 -8
rect 148 -42 306 -8
rect 340 -42 498 -8
rect 532 -42 690 -8
rect 724 -42 882 -8
rect 916 -42 1074 -8
rect 1108 -42 1266 -8
rect 1300 -42 1458 -8
rect 1492 -42 1508 -8
<< viali >>
rect 114 2322 148 2356
rect 306 2322 340 2356
rect 498 2322 532 2356
rect 690 2322 724 2356
rect 882 2322 916 2356
rect 1074 2322 1108 2356
rect 1266 2322 1300 2356
rect 1458 2322 1492 2356
rect 18 1812 52 1846
rect 210 1812 244 1846
rect 402 1812 436 1846
rect 594 1812 628 1846
rect 786 1812 820 1846
rect 978 1812 1012 1846
rect 1170 1812 1204 1846
rect 1362 1812 1396 1846
rect 18 1704 52 1738
rect 210 1704 244 1738
rect 402 1704 436 1738
rect 594 1704 628 1738
rect 786 1704 820 1738
rect 978 1704 1012 1738
rect 1170 1704 1204 1738
rect 1362 1704 1396 1738
rect 114 1194 148 1228
rect 306 1194 340 1228
rect 498 1194 532 1228
rect 690 1194 724 1228
rect 882 1194 916 1228
rect 1074 1194 1108 1228
rect 1266 1194 1300 1228
rect 1458 1194 1492 1228
rect 114 1086 148 1120
rect 306 1086 340 1120
rect 498 1086 532 1120
rect 690 1086 724 1120
rect 882 1086 916 1120
rect 1074 1086 1108 1120
rect 1266 1086 1300 1120
rect 1458 1086 1492 1120
rect 18 576 52 610
rect 210 576 244 610
rect 402 576 436 610
rect 594 576 628 610
rect 786 576 820 610
rect 978 576 1012 610
rect 1170 576 1204 610
rect 1362 576 1396 610
rect 18 468 52 502
rect 210 468 244 502
rect 402 468 436 502
rect 594 468 628 502
rect 786 468 820 502
rect 978 468 1012 502
rect 1170 468 1204 502
rect 1362 468 1396 502
rect 114 -42 148 -8
rect 306 -42 340 -8
rect 498 -42 532 -8
rect 690 -42 724 -8
rect 882 -42 916 -8
rect 1074 -42 1108 -8
rect 1266 -42 1300 -8
rect 1458 -42 1492 -8
<< metal1 >>
rect 2 2356 1508 2362
rect 2 2322 114 2356
rect 148 2322 306 2356
rect 340 2322 498 2356
rect 532 2322 690 2356
rect 724 2322 882 2356
rect 916 2322 1074 2356
rect 1108 2322 1266 2356
rect 1300 2322 1458 2356
rect 1492 2322 1508 2356
rect 2 2316 1508 2322
rect 2 1846 1508 1852
rect 2 1812 18 1846
rect 52 1812 210 1846
rect 244 1812 402 1846
rect 436 1812 594 1846
rect 628 1812 786 1846
rect 820 1812 978 1846
rect 1012 1812 1170 1846
rect 1204 1812 1362 1846
rect 1396 1812 1508 1846
rect 2 1806 1508 1812
rect 2 1738 1508 1744
rect 2 1704 18 1738
rect 52 1704 210 1738
rect 244 1704 402 1738
rect 436 1704 594 1738
rect 628 1704 786 1738
rect 820 1704 978 1738
rect 1012 1704 1170 1738
rect 1204 1704 1362 1738
rect 1396 1704 1508 1738
rect 2 1698 1508 1704
rect 2 1228 1508 1234
rect 2 1194 114 1228
rect 148 1194 306 1228
rect 340 1194 498 1228
rect 532 1194 690 1228
rect 724 1194 882 1228
rect 916 1194 1074 1228
rect 1108 1194 1266 1228
rect 1300 1194 1458 1228
rect 1492 1194 1508 1228
rect 2 1188 1508 1194
rect 2 1120 1508 1126
rect 2 1086 114 1120
rect 148 1086 306 1120
rect 340 1086 498 1120
rect 532 1086 690 1120
rect 724 1086 882 1120
rect 916 1086 1074 1120
rect 1108 1086 1266 1120
rect 1300 1086 1458 1120
rect 1492 1086 1508 1120
rect 2 1080 1508 1086
rect 2 610 1508 616
rect 2 576 18 610
rect 52 576 210 610
rect 244 576 402 610
rect 436 576 594 610
rect 628 576 786 610
rect 820 576 978 610
rect 1012 576 1170 610
rect 1204 576 1362 610
rect 1396 576 1508 610
rect 2 570 1508 576
rect 2 502 1508 508
rect 2 468 18 502
rect 52 468 210 502
rect 244 468 402 502
rect 436 468 594 502
rect 628 468 786 502
rect 820 468 978 502
rect 1012 468 1170 502
rect 1204 468 1362 502
rect 1396 468 1508 502
rect 2 462 1508 468
rect 2 -8 1508 -2
rect 2 -42 114 -8
rect 148 -42 306 -8
rect 340 -42 498 -8
rect 532 -42 690 -8
rect 724 -42 882 -8
rect 916 -42 1074 -8
rect 1108 -42 1266 -8
rect 1300 -42 1458 -8
rect 1492 -42 1508 -8
rect 2 -48 1508 -42
use sky130_fd_pr__nfet_01v8_A574RZ  sky130_fd_pr__nfet_01v8_A574RZ_0
timestamp 1646921651
transform 1 0 1251 0 1 -2767
box -1431 -2573 1431 2573
use sky130_fd_pr__nfet_01v8_ED72KE  sky130_fd_pr__nfet_01v8_ED72KE_0
timestamp 1646921651
transform 1 0 755 0 1 1157
box -935 -1337 935 1337
<< end >>
