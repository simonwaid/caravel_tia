magic
tech sky130A
magscale 1 2
timestamp 1645633816
<< pwell >>
rect -1457 -1119 1457 1119
<< nmoslvt >>
rect -1261 109 -1061 909
rect -1003 109 -803 909
rect -745 109 -545 909
rect -487 109 -287 909
rect -229 109 -29 909
rect 29 109 229 909
rect 287 109 487 909
rect 545 109 745 909
rect 803 109 1003 909
rect 1061 109 1261 909
rect -1261 -909 -1061 -109
rect -1003 -909 -803 -109
rect -745 -909 -545 -109
rect -487 -909 -287 -109
rect -229 -909 -29 -109
rect 29 -909 229 -109
rect 287 -909 487 -109
rect 545 -909 745 -109
rect 803 -909 1003 -109
rect 1061 -909 1261 -109
<< ndiff >>
rect -1319 897 -1261 909
rect -1319 121 -1307 897
rect -1273 121 -1261 897
rect -1319 109 -1261 121
rect -1061 897 -1003 909
rect -1061 121 -1049 897
rect -1015 121 -1003 897
rect -1061 109 -1003 121
rect -803 897 -745 909
rect -803 121 -791 897
rect -757 121 -745 897
rect -803 109 -745 121
rect -545 897 -487 909
rect -545 121 -533 897
rect -499 121 -487 897
rect -545 109 -487 121
rect -287 897 -229 909
rect -287 121 -275 897
rect -241 121 -229 897
rect -287 109 -229 121
rect -29 897 29 909
rect -29 121 -17 897
rect 17 121 29 897
rect -29 109 29 121
rect 229 897 287 909
rect 229 121 241 897
rect 275 121 287 897
rect 229 109 287 121
rect 487 897 545 909
rect 487 121 499 897
rect 533 121 545 897
rect 487 109 545 121
rect 745 897 803 909
rect 745 121 757 897
rect 791 121 803 897
rect 745 109 803 121
rect 1003 897 1061 909
rect 1003 121 1015 897
rect 1049 121 1061 897
rect 1003 109 1061 121
rect 1261 897 1319 909
rect 1261 121 1273 897
rect 1307 121 1319 897
rect 1261 109 1319 121
rect -1319 -121 -1261 -109
rect -1319 -897 -1307 -121
rect -1273 -897 -1261 -121
rect -1319 -909 -1261 -897
rect -1061 -121 -1003 -109
rect -1061 -897 -1049 -121
rect -1015 -897 -1003 -121
rect -1061 -909 -1003 -897
rect -803 -121 -745 -109
rect -803 -897 -791 -121
rect -757 -897 -745 -121
rect -803 -909 -745 -897
rect -545 -121 -487 -109
rect -545 -897 -533 -121
rect -499 -897 -487 -121
rect -545 -909 -487 -897
rect -287 -121 -229 -109
rect -287 -897 -275 -121
rect -241 -897 -229 -121
rect -287 -909 -229 -897
rect -29 -121 29 -109
rect -29 -897 -17 -121
rect 17 -897 29 -121
rect -29 -909 29 -897
rect 229 -121 287 -109
rect 229 -897 241 -121
rect 275 -897 287 -121
rect 229 -909 287 -897
rect 487 -121 545 -109
rect 487 -897 499 -121
rect 533 -897 545 -121
rect 487 -909 545 -897
rect 745 -121 803 -109
rect 745 -897 757 -121
rect 791 -897 803 -121
rect 745 -909 803 -897
rect 1003 -121 1061 -109
rect 1003 -897 1015 -121
rect 1049 -897 1061 -121
rect 1003 -909 1061 -897
rect 1261 -121 1319 -109
rect 1261 -897 1273 -121
rect 1307 -897 1319 -121
rect 1261 -909 1319 -897
<< ndiffc >>
rect -1307 121 -1273 897
rect -1049 121 -1015 897
rect -791 121 -757 897
rect -533 121 -499 897
rect -275 121 -241 897
rect -17 121 17 897
rect 241 121 275 897
rect 499 121 533 897
rect 757 121 791 897
rect 1015 121 1049 897
rect 1273 121 1307 897
rect -1307 -897 -1273 -121
rect -1049 -897 -1015 -121
rect -791 -897 -757 -121
rect -533 -897 -499 -121
rect -275 -897 -241 -121
rect -17 -897 17 -121
rect 241 -897 275 -121
rect 499 -897 533 -121
rect 757 -897 791 -121
rect 1015 -897 1049 -121
rect 1273 -897 1307 -121
<< psubdiff >>
rect -1421 1049 -1325 1083
rect 1325 1049 1421 1083
rect -1421 987 -1387 1049
rect 1387 987 1421 1049
rect -1421 -1049 -1387 -987
rect 1387 -1049 1421 -987
rect -1421 -1083 -1325 -1049
rect 1325 -1083 1421 -1049
<< psubdiffcont >>
rect -1325 1049 1325 1083
rect -1421 -987 -1387 987
rect 1387 -987 1421 987
rect -1325 -1083 1325 -1049
<< poly >>
rect -1261 981 -1061 997
rect -1261 947 -1245 981
rect -1077 947 -1061 981
rect -1261 909 -1061 947
rect -1003 981 -803 997
rect -1003 947 -987 981
rect -819 947 -803 981
rect -1003 909 -803 947
rect -745 981 -545 997
rect -745 947 -729 981
rect -561 947 -545 981
rect -745 909 -545 947
rect -487 981 -287 997
rect -487 947 -471 981
rect -303 947 -287 981
rect -487 909 -287 947
rect -229 981 -29 997
rect -229 947 -213 981
rect -45 947 -29 981
rect -229 909 -29 947
rect 29 981 229 997
rect 29 947 45 981
rect 213 947 229 981
rect 29 909 229 947
rect 287 981 487 997
rect 287 947 303 981
rect 471 947 487 981
rect 287 909 487 947
rect 545 981 745 997
rect 545 947 561 981
rect 729 947 745 981
rect 545 909 745 947
rect 803 981 1003 997
rect 803 947 819 981
rect 987 947 1003 981
rect 803 909 1003 947
rect 1061 981 1261 997
rect 1061 947 1077 981
rect 1245 947 1261 981
rect 1061 909 1261 947
rect -1261 71 -1061 109
rect -1261 37 -1245 71
rect -1077 37 -1061 71
rect -1261 21 -1061 37
rect -1003 71 -803 109
rect -1003 37 -987 71
rect -819 37 -803 71
rect -1003 21 -803 37
rect -745 71 -545 109
rect -745 37 -729 71
rect -561 37 -545 71
rect -745 21 -545 37
rect -487 71 -287 109
rect -487 37 -471 71
rect -303 37 -287 71
rect -487 21 -287 37
rect -229 71 -29 109
rect -229 37 -213 71
rect -45 37 -29 71
rect -229 21 -29 37
rect 29 71 229 109
rect 29 37 45 71
rect 213 37 229 71
rect 29 21 229 37
rect 287 71 487 109
rect 287 37 303 71
rect 471 37 487 71
rect 287 21 487 37
rect 545 71 745 109
rect 545 37 561 71
rect 729 37 745 71
rect 545 21 745 37
rect 803 71 1003 109
rect 803 37 819 71
rect 987 37 1003 71
rect 803 21 1003 37
rect 1061 71 1261 109
rect 1061 37 1077 71
rect 1245 37 1261 71
rect 1061 21 1261 37
rect -1261 -37 -1061 -21
rect -1261 -71 -1245 -37
rect -1077 -71 -1061 -37
rect -1261 -109 -1061 -71
rect -1003 -37 -803 -21
rect -1003 -71 -987 -37
rect -819 -71 -803 -37
rect -1003 -109 -803 -71
rect -745 -37 -545 -21
rect -745 -71 -729 -37
rect -561 -71 -545 -37
rect -745 -109 -545 -71
rect -487 -37 -287 -21
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -487 -109 -287 -71
rect -229 -37 -29 -21
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect -229 -109 -29 -71
rect 29 -37 229 -21
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 29 -109 229 -71
rect 287 -37 487 -21
rect 287 -71 303 -37
rect 471 -71 487 -37
rect 287 -109 487 -71
rect 545 -37 745 -21
rect 545 -71 561 -37
rect 729 -71 745 -37
rect 545 -109 745 -71
rect 803 -37 1003 -21
rect 803 -71 819 -37
rect 987 -71 1003 -37
rect 803 -109 1003 -71
rect 1061 -37 1261 -21
rect 1061 -71 1077 -37
rect 1245 -71 1261 -37
rect 1061 -109 1261 -71
rect -1261 -947 -1061 -909
rect -1261 -981 -1245 -947
rect -1077 -981 -1061 -947
rect -1261 -997 -1061 -981
rect -1003 -947 -803 -909
rect -1003 -981 -987 -947
rect -819 -981 -803 -947
rect -1003 -997 -803 -981
rect -745 -947 -545 -909
rect -745 -981 -729 -947
rect -561 -981 -545 -947
rect -745 -997 -545 -981
rect -487 -947 -287 -909
rect -487 -981 -471 -947
rect -303 -981 -287 -947
rect -487 -997 -287 -981
rect -229 -947 -29 -909
rect -229 -981 -213 -947
rect -45 -981 -29 -947
rect -229 -997 -29 -981
rect 29 -947 229 -909
rect 29 -981 45 -947
rect 213 -981 229 -947
rect 29 -997 229 -981
rect 287 -947 487 -909
rect 287 -981 303 -947
rect 471 -981 487 -947
rect 287 -997 487 -981
rect 545 -947 745 -909
rect 545 -981 561 -947
rect 729 -981 745 -947
rect 545 -997 745 -981
rect 803 -947 1003 -909
rect 803 -981 819 -947
rect 987 -981 1003 -947
rect 803 -997 1003 -981
rect 1061 -947 1261 -909
rect 1061 -981 1077 -947
rect 1245 -981 1261 -947
rect 1061 -997 1261 -981
<< polycont >>
rect -1245 947 -1077 981
rect -987 947 -819 981
rect -729 947 -561 981
rect -471 947 -303 981
rect -213 947 -45 981
rect 45 947 213 981
rect 303 947 471 981
rect 561 947 729 981
rect 819 947 987 981
rect 1077 947 1245 981
rect -1245 37 -1077 71
rect -987 37 -819 71
rect -729 37 -561 71
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect 561 37 729 71
rect 819 37 987 71
rect 1077 37 1245 71
rect -1245 -71 -1077 -37
rect -987 -71 -819 -37
rect -729 -71 -561 -37
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect 561 -71 729 -37
rect 819 -71 987 -37
rect 1077 -71 1245 -37
rect -1245 -981 -1077 -947
rect -987 -981 -819 -947
rect -729 -981 -561 -947
rect -471 -981 -303 -947
rect -213 -981 -45 -947
rect 45 -981 213 -947
rect 303 -981 471 -947
rect 561 -981 729 -947
rect 819 -981 987 -947
rect 1077 -981 1245 -947
<< locali >>
rect -1421 1049 -1325 1083
rect 1325 1049 1421 1083
rect -1421 987 -1387 1049
rect 1387 987 1421 1049
rect -1261 947 -1245 981
rect -1077 947 -1061 981
rect -1003 947 -987 981
rect -819 947 -803 981
rect -745 947 -729 981
rect -561 947 -545 981
rect -487 947 -471 981
rect -303 947 -287 981
rect -229 947 -213 981
rect -45 947 -29 981
rect 29 947 45 981
rect 213 947 229 981
rect 287 947 303 981
rect 471 947 487 981
rect 545 947 561 981
rect 729 947 745 981
rect 803 947 819 981
rect 987 947 1003 981
rect 1061 947 1077 981
rect 1245 947 1261 981
rect -1307 897 -1273 913
rect -1307 105 -1273 121
rect -1049 897 -1015 913
rect -1049 105 -1015 121
rect -791 897 -757 913
rect -791 105 -757 121
rect -533 897 -499 913
rect -533 105 -499 121
rect -275 897 -241 913
rect -275 105 -241 121
rect -17 897 17 913
rect -17 105 17 121
rect 241 897 275 913
rect 241 105 275 121
rect 499 897 533 913
rect 499 105 533 121
rect 757 897 791 913
rect 757 105 791 121
rect 1015 897 1049 913
rect 1015 105 1049 121
rect 1273 897 1307 913
rect 1273 105 1307 121
rect -1261 37 -1245 71
rect -1077 37 -1061 71
rect -1003 37 -987 71
rect -819 37 -803 71
rect -745 37 -729 71
rect -561 37 -545 71
rect -487 37 -471 71
rect -303 37 -287 71
rect -229 37 -213 71
rect -45 37 -29 71
rect 29 37 45 71
rect 213 37 229 71
rect 287 37 303 71
rect 471 37 487 71
rect 545 37 561 71
rect 729 37 745 71
rect 803 37 819 71
rect 987 37 1003 71
rect 1061 37 1077 71
rect 1245 37 1261 71
rect -1261 -71 -1245 -37
rect -1077 -71 -1061 -37
rect -1003 -71 -987 -37
rect -819 -71 -803 -37
rect -745 -71 -729 -37
rect -561 -71 -545 -37
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 287 -71 303 -37
rect 471 -71 487 -37
rect 545 -71 561 -37
rect 729 -71 745 -37
rect 803 -71 819 -37
rect 987 -71 1003 -37
rect 1061 -71 1077 -37
rect 1245 -71 1261 -37
rect -1307 -121 -1273 -105
rect -1307 -913 -1273 -897
rect -1049 -121 -1015 -105
rect -1049 -913 -1015 -897
rect -791 -121 -757 -105
rect -791 -913 -757 -897
rect -533 -121 -499 -105
rect -533 -913 -499 -897
rect -275 -121 -241 -105
rect -275 -913 -241 -897
rect -17 -121 17 -105
rect -17 -913 17 -897
rect 241 -121 275 -105
rect 241 -913 275 -897
rect 499 -121 533 -105
rect 499 -913 533 -897
rect 757 -121 791 -105
rect 757 -913 791 -897
rect 1015 -121 1049 -105
rect 1015 -913 1049 -897
rect 1273 -121 1307 -105
rect 1273 -913 1307 -897
rect -1261 -981 -1245 -947
rect -1077 -981 -1061 -947
rect -1003 -981 -987 -947
rect -819 -981 -803 -947
rect -745 -981 -729 -947
rect -561 -981 -545 -947
rect -487 -981 -471 -947
rect -303 -981 -287 -947
rect -229 -981 -213 -947
rect -45 -981 -29 -947
rect 29 -981 45 -947
rect 213 -981 229 -947
rect 287 -981 303 -947
rect 471 -981 487 -947
rect 545 -981 561 -947
rect 729 -981 745 -947
rect 803 -981 819 -947
rect 987 -981 1003 -947
rect 1061 -981 1077 -947
rect 1245 -981 1261 -947
rect -1421 -1049 -1387 -987
rect 1387 -1049 1421 -987
rect -1421 -1083 -1325 -1049
rect 1325 -1083 1421 -1049
<< viali >>
rect -1245 947 -1077 981
rect -987 947 -819 981
rect -729 947 -561 981
rect -471 947 -303 981
rect -213 947 -45 981
rect 45 947 213 981
rect 303 947 471 981
rect 561 947 729 981
rect 819 947 987 981
rect 1077 947 1245 981
rect -1307 121 -1273 897
rect -1049 121 -1015 897
rect -791 121 -757 897
rect -533 121 -499 897
rect -275 121 -241 897
rect -17 121 17 897
rect 241 121 275 897
rect 499 121 533 897
rect 757 121 791 897
rect 1015 121 1049 897
rect 1273 121 1307 897
rect -1245 37 -1077 71
rect -987 37 -819 71
rect -729 37 -561 71
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect 561 37 729 71
rect 819 37 987 71
rect 1077 37 1245 71
rect -1245 -71 -1077 -37
rect -987 -71 -819 -37
rect -729 -71 -561 -37
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect 561 -71 729 -37
rect 819 -71 987 -37
rect 1077 -71 1245 -37
rect -1307 -897 -1273 -121
rect -1049 -897 -1015 -121
rect -791 -897 -757 -121
rect -533 -897 -499 -121
rect -275 -897 -241 -121
rect -17 -897 17 -121
rect 241 -897 275 -121
rect 499 -897 533 -121
rect 757 -897 791 -121
rect 1015 -897 1049 -121
rect 1273 -897 1307 -121
rect -1245 -981 -1077 -947
rect -987 -981 -819 -947
rect -729 -981 -561 -947
rect -471 -981 -303 -947
rect -213 -981 -45 -947
rect 45 -981 213 -947
rect 303 -981 471 -947
rect 561 -981 729 -947
rect 819 -981 987 -947
rect 1077 -981 1245 -947
<< metal1 >>
rect -1257 981 -1065 987
rect -1257 947 -1245 981
rect -1077 947 -1065 981
rect -1257 941 -1065 947
rect -999 981 -807 987
rect -999 947 -987 981
rect -819 947 -807 981
rect -999 941 -807 947
rect -741 981 -549 987
rect -741 947 -729 981
rect -561 947 -549 981
rect -741 941 -549 947
rect -483 981 -291 987
rect -483 947 -471 981
rect -303 947 -291 981
rect -483 941 -291 947
rect -225 981 -33 987
rect -225 947 -213 981
rect -45 947 -33 981
rect -225 941 -33 947
rect 33 981 225 987
rect 33 947 45 981
rect 213 947 225 981
rect 33 941 225 947
rect 291 981 483 987
rect 291 947 303 981
rect 471 947 483 981
rect 291 941 483 947
rect 549 981 741 987
rect 549 947 561 981
rect 729 947 741 981
rect 549 941 741 947
rect 807 981 999 987
rect 807 947 819 981
rect 987 947 999 981
rect 807 941 999 947
rect 1065 981 1257 987
rect 1065 947 1077 981
rect 1245 947 1257 981
rect 1065 941 1257 947
rect -1313 897 -1267 909
rect -1313 121 -1307 897
rect -1273 121 -1267 897
rect -1313 109 -1267 121
rect -1055 897 -1009 909
rect -1055 121 -1049 897
rect -1015 121 -1009 897
rect -1055 109 -1009 121
rect -797 897 -751 909
rect -797 121 -791 897
rect -757 121 -751 897
rect -797 109 -751 121
rect -539 897 -493 909
rect -539 121 -533 897
rect -499 121 -493 897
rect -539 109 -493 121
rect -281 897 -235 909
rect -281 121 -275 897
rect -241 121 -235 897
rect -281 109 -235 121
rect -23 897 23 909
rect -23 121 -17 897
rect 17 121 23 897
rect -23 109 23 121
rect 235 897 281 909
rect 235 121 241 897
rect 275 121 281 897
rect 235 109 281 121
rect 493 897 539 909
rect 493 121 499 897
rect 533 121 539 897
rect 493 109 539 121
rect 751 897 797 909
rect 751 121 757 897
rect 791 121 797 897
rect 751 109 797 121
rect 1009 897 1055 909
rect 1009 121 1015 897
rect 1049 121 1055 897
rect 1009 109 1055 121
rect 1267 897 1313 909
rect 1267 121 1273 897
rect 1307 121 1313 897
rect 1267 109 1313 121
rect -1257 71 -1065 77
rect -1257 37 -1245 71
rect -1077 37 -1065 71
rect -1257 31 -1065 37
rect -999 71 -807 77
rect -999 37 -987 71
rect -819 37 -807 71
rect -999 31 -807 37
rect -741 71 -549 77
rect -741 37 -729 71
rect -561 37 -549 71
rect -741 31 -549 37
rect -483 71 -291 77
rect -483 37 -471 71
rect -303 37 -291 71
rect -483 31 -291 37
rect -225 71 -33 77
rect -225 37 -213 71
rect -45 37 -33 71
rect -225 31 -33 37
rect 33 71 225 77
rect 33 37 45 71
rect 213 37 225 71
rect 33 31 225 37
rect 291 71 483 77
rect 291 37 303 71
rect 471 37 483 71
rect 291 31 483 37
rect 549 71 741 77
rect 549 37 561 71
rect 729 37 741 71
rect 549 31 741 37
rect 807 71 999 77
rect 807 37 819 71
rect 987 37 999 71
rect 807 31 999 37
rect 1065 71 1257 77
rect 1065 37 1077 71
rect 1245 37 1257 71
rect 1065 31 1257 37
rect -1257 -37 -1065 -31
rect -1257 -71 -1245 -37
rect -1077 -71 -1065 -37
rect -1257 -77 -1065 -71
rect -999 -37 -807 -31
rect -999 -71 -987 -37
rect -819 -71 -807 -37
rect -999 -77 -807 -71
rect -741 -37 -549 -31
rect -741 -71 -729 -37
rect -561 -71 -549 -37
rect -741 -77 -549 -71
rect -483 -37 -291 -31
rect -483 -71 -471 -37
rect -303 -71 -291 -37
rect -483 -77 -291 -71
rect -225 -37 -33 -31
rect -225 -71 -213 -37
rect -45 -71 -33 -37
rect -225 -77 -33 -71
rect 33 -37 225 -31
rect 33 -71 45 -37
rect 213 -71 225 -37
rect 33 -77 225 -71
rect 291 -37 483 -31
rect 291 -71 303 -37
rect 471 -71 483 -37
rect 291 -77 483 -71
rect 549 -37 741 -31
rect 549 -71 561 -37
rect 729 -71 741 -37
rect 549 -77 741 -71
rect 807 -37 999 -31
rect 807 -71 819 -37
rect 987 -71 999 -37
rect 807 -77 999 -71
rect 1065 -37 1257 -31
rect 1065 -71 1077 -37
rect 1245 -71 1257 -37
rect 1065 -77 1257 -71
rect -1313 -121 -1267 -109
rect -1313 -897 -1307 -121
rect -1273 -897 -1267 -121
rect -1313 -909 -1267 -897
rect -1055 -121 -1009 -109
rect -1055 -897 -1049 -121
rect -1015 -897 -1009 -121
rect -1055 -909 -1009 -897
rect -797 -121 -751 -109
rect -797 -897 -791 -121
rect -757 -897 -751 -121
rect -797 -909 -751 -897
rect -539 -121 -493 -109
rect -539 -897 -533 -121
rect -499 -897 -493 -121
rect -539 -909 -493 -897
rect -281 -121 -235 -109
rect -281 -897 -275 -121
rect -241 -897 -235 -121
rect -281 -909 -235 -897
rect -23 -121 23 -109
rect -23 -897 -17 -121
rect 17 -897 23 -121
rect -23 -909 23 -897
rect 235 -121 281 -109
rect 235 -897 241 -121
rect 275 -897 281 -121
rect 235 -909 281 -897
rect 493 -121 539 -109
rect 493 -897 499 -121
rect 533 -897 539 -121
rect 493 -909 539 -897
rect 751 -121 797 -109
rect 751 -897 757 -121
rect 791 -897 797 -121
rect 751 -909 797 -897
rect 1009 -121 1055 -109
rect 1009 -897 1015 -121
rect 1049 -897 1055 -121
rect 1009 -909 1055 -897
rect 1267 -121 1313 -109
rect 1267 -897 1273 -121
rect 1307 -897 1313 -121
rect 1267 -909 1313 -897
rect -1257 -947 -1065 -941
rect -1257 -981 -1245 -947
rect -1077 -981 -1065 -947
rect -1257 -987 -1065 -981
rect -999 -947 -807 -941
rect -999 -981 -987 -947
rect -819 -981 -807 -947
rect -999 -987 -807 -981
rect -741 -947 -549 -941
rect -741 -981 -729 -947
rect -561 -981 -549 -947
rect -741 -987 -549 -981
rect -483 -947 -291 -941
rect -483 -981 -471 -947
rect -303 -981 -291 -947
rect -483 -987 -291 -981
rect -225 -947 -33 -941
rect -225 -981 -213 -947
rect -45 -981 -33 -947
rect -225 -987 -33 -981
rect 33 -947 225 -941
rect 33 -981 45 -947
rect 213 -981 225 -947
rect 33 -987 225 -981
rect 291 -947 483 -941
rect 291 -981 303 -947
rect 471 -981 483 -947
rect 291 -987 483 -981
rect 549 -947 741 -941
rect 549 -981 561 -947
rect 729 -981 741 -947
rect 549 -987 741 -981
rect 807 -947 999 -941
rect 807 -981 819 -947
rect 987 -981 999 -947
rect 807 -987 999 -981
rect 1065 -947 1257 -941
rect 1065 -981 1077 -947
rect 1245 -981 1257 -947
rect 1065 -987 1257 -981
<< properties >>
string FIXED_BBOX -1404 -1066 1404 1066
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 4 l 1 m 2 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
